XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
N�'��`�'ɽ(�\b4��[6���\M��Ţ���8P�xI����!� p�fT&�8��~�N��)"��;۠Z$����z>e�C�އ�A نq�A�H��4�Μk�?��;������8c�W������&����#7WJ(��@�*�:�o%���<��&���	�IyL��j��ע�G�Nh�ӕE���ɛ�Ġ�ve�?����G ����g;^�r�Ŕ>���?��Π&�xojs�qR�).킽!��M;�x�_����G`�nbt�U�"��}C8G�x���"�hڇ�5������Q��Z�5��Vf�LF�d���-6}L~�m�����L��+Q�y�߼���^KϬ�lF^A�47���p�c��E{?��ɵ�J�_�O���k��-Sx'��L%À�٪I*�D�S��S�e���{	�&W+�	���i������0�����g�n�����ett�#|��JhR�N���٭�R��M4�SB�+T��� 6g9��ޤ�
��$S�1,]�,FqNB�n���r1�c� �70L_2F+b��I�U���p#�e�e�9������e[�SP�������֥�nX��{;EX{�|���5;6�L�w5�2�Aq�;!��������K�I�ՈX5���+��'�h��H.�W��?QP���G���m~Z����l!��:���d��������ɕ�r	�q�o����8�����Αg�H����Ɲ�Zo��(�XlxVHYEB     f6d     6f0E�	R��P#���=�b�L��|�荊��v�^a%�������xj~K�T",W�8���φ��a���������'#�J���!�y��.�gC�cD���|U��G`���G|��^��h}�N�N4ձ��>�jq������?F3kZ�Q��6hA�Ҏ*�%�\��NEma�C��l��]X��i]0��q��Z
X�SY���/������%e��ϩ2�z�cYz`AHj��>�������G矙�2�R��Z�Sn��g�7m��vn͉�
��X�@7M���8kch�=PKv.1:8B�f�t�{���04�X'�>�y�@��Ӆ6�~ԝ5i{pB����	V��������E5D�o�*�����.#�<�7�ά���e�4Y؝O,���\f5�>�y��.*�@�^%�9B�Ccl�3¹zL�^=�q6��0az�B�gU;��zn#�ɼ<��Kt�<������_���ẘ!����s�4�5n��	~j]B��E�ԋ	�
+��|`��X�`�&:єa���K��7;�N�c5)՝׸b6'�����60�X� ��w����$ĶC��*љ�2�Mq��F2�"uk��`�.P�f6������ �۹��h�n��K��Q]��-q��)6�X�U�<c[�G3�|&����&
�3d�1
ّW�r�aP�=��~������(���$[�Ш8m�U2�M���k=��,��{hݰ�l�#��8<̛?q��WuqCq&�q�H��Г�\���B,��7����"��ij?
{�X���k����a2�>�OC7��!������f�'�oՄ��E��&b�Qqn㇀��QbznPm�W{2�
�B��7�H;��Ȗ�~CXqK\���fX�98�V��hCn�Ey�S<����\g8��R���:䇪}Y�-usD��_~n���t��������#���p�WYjDY�n#N�ge�NWe!K����BHV�C~�'��r#"�����G�w��C�{�� �J�'H�}i��ؖ��۸�U�`X�m�m�p��(��@�[u_�}?�3�b�j��K	�k���n�K����5�]�YX1R`�*ɬR����$�S	��(6�Y�X[��V���X\=
ȫn�xORes�7�x����>�x���3�?\٩��p�'�-����!�Iv���I��H8�4��,�Cb�"�����p_'�be(c�aT�b�����b�G �(�Nh�%��4}���(8Y�y�G���>�kL�ǋ�.��A��`�l��������ۤ���8ƃ���ԙ�!xV �`�����
goX粪!Fu88/b'eŝ\.)�ǣ�@3�ߦ��V8e\�%#!�؛צ�kL(��<�d0j�@[Ȗpb�ߎ
���c
��q���>�͖��:���������l�.�-�Bo�^�S��#�1�"�!mWu��Wy,�4�2� `>����_~��;�{KݢX b�ю�M�G��ZbƄ8쐨��֚�w��fӪ�J��3q�{;��;ƞ����\]��q�6t�0��-��t!q��e�besi��d�����3����_����RL7�|1�N���޸6��&|'{n�_��1�.a~J�Я<`}ԯ͈��}�S�Ѡ�s���S�Gc�^�(+$ �IL�
vH��̩�*����7@E�����P*��0���1Qq�Tǻ ����}��/O��з��