XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`H������~��d�e2��ݳAM�hCZ]�푍R%ҳ'0Le�e�!�ki�-�k�V��^���a��(�S�{J�T)�^5gU'9��$����yi53le�V�� s*�_z���!:�~�8�B�wg1��A�'m�m0�wQ3k�����|(g��#ꡧL�U�@E9`��@��b�(N�#�+��'ao�^~8;� �lO�E]�f�P�}ޖ	�̨�M��T����>�afp |TO�l�=fŁ�ћ|�S�g��+x�­�ɷM�R�.��� �
u��L�����F�
08j���x�Z#%�j�!������<2�
��/qhY����ܘN�y���ʚ�������e��1h�J�R`�CDL��:�������J���u��t�̮%:�;��U²��( ��Ղa�R�k�o`0��LFް�Ƶ}�ع���]�T\� ���ꛫ�+��p�`$�
��6[,�-����1�j��DU�Px�ز���{���דQ�Ƅ��G����𿡒GJ�����9)��<̺��d��VA��T(�91ķ�9k�ƙ��s�K��CG�"/�kd�"�F�^�;;i =%�
��Lf�N�"�<_�{uM,l���ۼe�mE|����Gs������267A�hu�':��r7�Y��
�pD�&L����y�On��� ˸���*Շ
�C5��;u��7h��w	�Wq�.�/d�^�SUs�n����OJ��q;�Ud��*Rq�o.�T2y�K��y�SXlxVHYEB    a037    1fe0cک�fWy�tK�	b�?�C�sv�3���d��غ�,
�7FvF��z즅�%�S�J��D�.@{����&b!W�?��>̨"���{�������hF*�6���V��/Nߵb,�`�zTtG�厵�s����1����oNf窲.�H�'&AHp���hQ��Bu a����6ґ��s�5�0�TG������yS��W�b�K�	(;���)Eb���[9���!�>�?"o��#'�~V���q��i'̸�D���1�ͮ��@���Sx����-1�ߒt���Pw��3�`Aө�P�1��k�r7s�E�;�6�WquWn[v2��it����3p��.
���u�s���U2|uc�`/m���v�����7��Ƹul�*4p��^2��)Or��Tή�24�fIa|7�{Fr�"��P�(����'��D�l>yY�R�ы��h�%G*�O��㌒�ʈ�]��ȸ������oV�z3��Gxx.N����KHI=K%��k�ݔz���F��$��o�Z��2�]�Vr�� 0^E���gE�.�V_����� nM���!f'�~�-��t��*J��`��e��&	������ݖ�K���ʢP�E���cV/�i�bf�)a@��|r��bI�\�p E�����~e������mX�xIм�vu�\R��ǆ���4PS���0�q�g&ڋ~�0A>�wL�~�d��3:c���@N��aō�q�weK��Y������P�HD�+L�m�D���9hG�/V/ȥ��&	�pt�P΀������
_��Y�n �0m�WPҙ���nw	q{ዢ� ����ZJѼ}r�OK�� �.�� 8IҷlN�qe��ki&�k�$�=��}SNq�,�W���Ġ��fɃ�&��PwE��UP�v�B��xK�����:�Z�U�7ϖ�{�]�HZ|A&~Y ��r�[Y�0�@"��0ʀO����_'Ek�$��k��Am	����?�a��RL�����&�]%
��O T�
FhT�@/�A�-��@*)��s[�D��Ӣmn.�eNto��vP��j���j�ĩ�a!_+�u�,6�)`���b��eׂ�4%��&Ajb�8�t1��imK���XG�(�hT�G�Բ�o�ŧ�;�%����<7�g
�73���#`k�9�OɐD4Ԏ�R1,�,�"e�P��\��Ȑ�������W�[5k���A�fao:�a��]���#��7%�ܾ��yYL �R"
�zԖ [5�+�1y!^�
��֞YsL�� ��A�Z�jñ�^y���;��>�?G���ɭI-�
t"��}A�������\�/0* 4#~�d�uZa�x�wT�����[�KH��1�SF�T��V	c�y¿�b���gy���T��l�f�"���-�iЇP
����N�?&H�yw����K����x���U�Ps�2��*���i��v�6��Ǩ+�t
4��F ڬ�Z'D(��)��H��ߕ]hpk�c�����ʉ^���?��O^�$��C	� xy/;aQu��0�����`p˨�^��h������_^���Z f�ڶx�9b��j����m6����~����B,✎��C��6g�$���EX�۫B֎�eޭS"X�C�@,��'py5l�i����>X\�G�������N�]ǅ밍�*��V`�<D@bn⨡���orߓ������Rr�ݰ|�072����Wv�L�|�rÆ&���C)f_<��v������;7\ݤ=fܔ����TJ+��,e��ê +�o�Yګq���y+$���%�f����
�X���8�#�gD���X]~��+���=���>�J����m�]�h}�����U���1��]"� ��>�r�&��w�J��XQ-�}��jWD^%V��/y�1&pζ����a�%�.x���& ���p�SV[���H����V�吐nX�k�.�y3�Ӡ�����i�B��u4�H�71;�n{ѧ���|�s�������b��(�v>{Yn���j��I���j��Y�&�ȸ�6�Ɏ�ر��(T��K(]��&g��u�N8Y���q�������	�(�h�'<���7�`~���Z�'�����{�{�0!O\��!Q�F8'�-*^a�i# ���3İ����ȕ�[�$�6��>��r��qﳺo���$�۞~s��n�ù�C�E%���B��}I�GY��
�o����XC��V8VnI��pt]��ҽ/C���6/��ulK�C�;�
On��o�0��(Ʃ�i�v6rD���7�z���xd|	^��ʾц?
׷��^!/��j�\DKf>�p��M�}�Z§Ų�Q6�4��t]�����Q���F������1͇����qR��h	�*9I�T�J�ʐ�+1���<P��}3��V�kN��7
DQ�FV��'i)@8�
�a��J��"��)L�JDM�Nk<��������s��d���[Y�?��߇�\��pZ�1bN)��KF��ς���|�a��{��G��]"��~yI���=�ie��+�`(�|\"�Θ� َ����u������d���=K����\�d[��4�ߚáë䚣-�7z[��;���j�8ě�c�^O&�Tiu_�/P��7O�l�L�b����f�KrYdhC�t���_G��HH�Kv�6�s^��餈���t�l(��]�ԫL������|Ҧ͎��Vs���)��TG.ؘA�[�w�kl�2�:��ƞY��i  Y�kQ���|3�G�!�l�Eͅ.A\oL�s�{��Ա�<��.R.F-9˥�8ﵮ�G��6n�_<>�m���Σ)�C�BEl�����ص|c�!ߖԑ��hQifB'2�Z:ı��9.��}a��u^&��/���+��K)����)b����H:Ѐ&�s�yz���'xXMH�	b�Ӥ�O���tn��XН���[���E��������1��^�>��_X��<i�	h�}<���ד	&�;��Z�Zh �qV�	{�#O���}V��?�*�)I��j��ۤ�_�9���ZX.�����;��А�W�}����1֔ Z��#LG��]����'҉�d5�3� ���8.S]�䆍'*)=/$>����e���\=	��⋥<9���e��`.MJ�(�;�t��$��yS�c+�L���f���J�s��N���S�Lޑ�n"ƫZ^Q�F�*����J
��@��B����]�Q�� _8�f��u>��9�n�ֳM����-q���l�2Y�
ŗE��i6�L��po(�x� �&���� eFN��qĿ��Ճ�`F-wT���cP�Y���)��&����
u?�aw�U���di:g�6���z2rF2��:s|�Ѕ`R�-��"�<,�-$��i�C�첄�q�NҜ5�dECk��e\�n�eEB��	@~GT�0Z���p]��쪱U�0�5�4��(���pgV�,%(�5��s[�?P�2Bs�MZd��?G<U��d`⸑�;�~��%~���'�H��q�8�[�]^κ��k:���]���a��WDg-������#�x|_�H��aXd�id����݃�x����3L�]|e͝-�?�Ck@#��;<������3�M�^�&�����d�� <_՚}KC�lql�j�S-)]�ך��~�{Ҧ�@xK�x)�|}H�GZO�����L��g�N����po!so� �J�5&��y�>��ήb��B�*z�2��> )6��qO�I{^���������/��#N伹R��o��,<D��7�����/H��|��\F����A����m��8���qSNTxU%��uYd�����3:��I��
���B�)q�O4�H+%2�2ҫ����2�A�,ڟ���H�H����JߵKX*�S���,���$Q4�0?J�>�����;�R�	/��Ny)#w����f���x� 
w���5�9��A��eg�6o&�瀷M���a� ��5u���.��]����F�OY$M*�Z������-�F�G���`��Aن�%t�����Y�:G[Ƨo�Q�on���r���#j�~���l�O��AV��h;ԴpL��FP2e߯�BrrtK������
��d�R�a���2]����_|w$�����{�)����0/4�.I|L���l�?,S�J�K��OYm,Td�IV��6�3�(}뷀5�;	e#9a��B���Vy]�hݴu��y��`$�(�CL���������!s�PNYc�7~HL_�w�R̂Q�@/�/�=%�P�2X}8'B�T��S� ��Cƒ�:�v���DNS �
%�� ��rT6�V��K{�l���ؒr~����D�� �EF\���1W�X�A��̠�YEIKTS�3��'EZ$�=�Z3�J��N�Qi�v�}󃎹₭���Qf7�M߹�>4~.�՝�����H�����[N��� ���������u�d�#�4�J6^74�^�b#&���BN�.�-J"*�i+({tc&KQ��%BQ6�Z$L�s��`�>�6r�;�{��fpU܀���ظ���c[�B�̔�Y4�n&&%��J؜e%][�B^e;۷\4{�w ̸���YS��Ц��K�b�o�ލ�J��Xr<�/hS�7��8��E(��Q/���5،F:�ȇU��'�\P�#R�V[��m�\YfH��e�j�@'�"���G��Z�N�c�7���=D�̹I~o���Eo��M��7s��نZpN�q�<-����4E)Y����8<��^�-���͞$���޵���~���Kmt���������l$�cJ3��':�G(�7�E���S���1o~�~���`<F���`��[����{�2h#P�B�T�[���:����I��d }�f�����{'v9"�e�R;�[�4������۾�y�ŝ������zܨ�{�\�f)�3/����z�Oρl)��c/whʡ�b�
޶���#�>��뛤:#�E�:��;"[���\ů�x05̹���#$Z����@�O{O�Ǟ��K:�`�C�v��Ҷѽ�MQ���n.��];C��O\�#����e���Ŋ��}���2�Y[��J�Y���RG��#�_@���=Tg㘉AGJ�t�.)��/��!�xTQ�X��\p�<��m�:!�Yp�� 䫵�M{�qr�p�N�R��/!��� �#�k;�3������%�<���m)�.�Ѯ�{��`Rr�$��7��cPf��+�'�6��9qN'�v��r^�1�[7��9�X�'��QyaD$�j�"a��V
��3�H��|,�0+�I�E^��i7�J��E�6�`��<Ef�Ύ@GEXwJ��(���=�5�����nј�{p�R���͊#5;�L���S�˩�)rX��KO2�����N�t� �,<0֝w�w�U�; �����$��v�������\��M�����(:K�&�r� �ys�א6s�zbƁ���J�d��>�ʘ��LJU��A0GZL�Ȋ�@�Xӳ��/O�3����8�l����T2�������e�N&*d<�)���2�HC��m��[l�>	�&�?�o\���%����5���i��2?P�Ȯ8'����a��9�z�W(f��t.݅Lֽ��v��j�pU��~�ʦ��A40���7�̻d��6>r�ߐÆ	~wSJF�A�/��3>����b2�nP ��{o[�Rf��g�ʙ2��-�q�j*�X��	}�n�LRy�׋�a�G)vz.��^�%�i��)�{V��=B�'F���\<�+���I#D��G� �։��!؆�A-����~8ɼ�%����@�t�k�^�y�J~�S������x��`��H>(�`@)^���̂*[T����Q��ẍCI.{K�x���r.����Q�% }"=�E^�M!OTK|�_�{�{��KE�C;E"'E�G��UiG�+����B�+X�S�]WX{A�W�C��̜��*wf'��l����j�����Bx#MΧC��?��/S:�!��]�o!�� ݱne4��?Cs�+|L2�"�=t�=������/y*ڔ�v�T��������=<����J{X ��!q��5�"�y����Ζ\m����z/4L`�����
��.��u{���0��v�(��g�
X�c�1�Lթȼ	�m��Y��	+X3������d�����Uf�!�`H�K�`G^<u�. �p�������1ݷ�oO8=H�=#��W�9k���d���2z-�y`�ᮊ��Xjq9� �\\?7�$)S�ꃖ^.:Ӄ+u���)@Bt��0�[?�j��"���#���E��C��d�\D�؍��G6��UD����n#Փм���0�_CH2��E���R}�¿Q	��nB{Ӽ�o���Uk�Hac�Rh`�1� �m����w�����K�E~������ )��J��u�V��G�傹�$�n]��`��>Ⱥ�j@S]�{� x�2l��ϐ������������߈V��6On�1�^���"�� �@ʵ���/�&�������2�b��^�V��+�e
�]'��	�9c��#�m�xcw���OF������h��n=gqi�Q�}�˻�H�=|hhtQ�����$�ӫ�4+4�Idt`�d�d�	�m��~j�ع�o�@�̿�Q¹�F�I��8��z����Zr��[��%{���[�zГQ�N����YEƨ|BQ���Ҽ&_�X�jn��{-��ɱ�r�����7�u�&J沲s��~�ld:$�	�oʦTcC�8�-�wlüln�d��m���x��Ag+H��XX^��-ٙS^���!���m�!�؊O����m�i �vi�qm���4�6�QZ'K�����rd �f��ƹ�q8��xX<�@�MN��y ���&;��ct�S�|�
,���S�}"���h� ��.�NV8���!S<�����
�z�4������9-�vy �'E�h;���F��a1@��q�v� ;��p"�<l��x��)']�.ERI(�I��a���FLj�R�HO\Jd4���@��j�m����&�j�?��ox��;����Ӳ��X�aK7��.JR���ޥ����,��݇W,��'�~�b�dV�E������9bi��<�k!���K��%pA:�ئ�7�C@nV$���� �d��C����&�&*T5����,��a�d�!Ӟ��pTE�,�>�}1�lĴ^>;Sm:\�qn�����E�R`��fA2�R/3�j[h('wd���^H���sm,թ���5$�ʕ=����1#���7d;H-]qӢY��EohӃq��x�`˂�103{R��T&������|�\���K���qy�.�2=���@�'�u6�)S @ �����CU0�f��b(5�`k���M�Y��:j�lHd������L�eW��� �y���Fq���* [��x�geW_��-�	��[��W�-*]�-fR���H�ÌI���9x8���!��}s�Cm&є�k�~�J� �I"�p�~+3ܺ>�B�m����[~r/A��
�=��.��O��v���uCE�!�GjM�5ٓU�/᧵��0�=\�W�P؞������S�c0�N�nOp����I���W���σ-Q��K�xГj�N�۲_�!`�/Խ{g2��&����S'SH��$aRT��N�R��sL�XLڢyf2{�����oHBu�f'^������]Ӧ������;�����[?&i��$w��H�|�W���bʆOqi�GJ��T���Q|f�1̣3֌�t�B�I+<�z������a2�Hu���6�%���3z���{}�[��0v��9��O�C���Y��ښ�UU%#R��}�6�.,7��������8�ښ]Z
D�	P
~�����t�Jv���mp�U@�[���Ц�yd��yn�ZH��"�Wz��\���