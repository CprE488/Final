XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ӹ���K�a����y-�ν]��]2�g���:��pC�J����f�*���0+��e���V�m�!�M��ť]��v�⚙�h��Cb�q��|1�H.�ڬ����B踡N�����,�%f�qFc0*X����+&J�*�ǰ�j�,J{��;o�����W�b}���Ho~�hm��^j+��'D��a�����N����4A�ܯ�Sk��)酢2�A����W4*�S(����Q4��b�5趟��V�����Z�瀨*�+�"�I]��J�F�����A���e�B.Y��)�ǩŚX���cט��R4�KM���I��
?+��D�uB���T����I�a�vwc�i�d�g��=q���R5���ŀ^�`�e%�Tm��­Q��5�qPˡJ���w�Fa!*��Y#\�#����M��H���� $�U��Q3��+����/u��d���'=2�T�d�±�G��C�k�w䭤�hX�&�mh����RA���ܬ�ʦM�a	��Qo�z�Bɬ!�[Јz��xa�bXK��B�ő����������H�'��YwM�Ŧq���5R����J3�*�E彩�R�G�h���?�7����V�],�UT�|��8vc������.�{B"����A�qT��~Bz��S��ͪ�~d�-�hV�E�hgFw��;��t�k��b����`�w�%&Rݲ�V�y�Zm�33�!�[Qda70�+��cJ��c��A:GmR�Qժ�q�XlxVHYEB    42ae    1110D���$p���H�=J�JE�틦��Ӽ��"�+��V���8䌹ɭ���I�^I�Z�17Cb�(l��W4�*�uˈ!+|w�8>�;��G>�q�+��\j8�Y�c��������t�j��|�i7�xú��K�>2�7��`�_��=c�O�ϭ)�꺃��3�|,�}S���,{G���n�]���g�歬^"�eTE���Ĺ�|��O�YG5�W�"z�0p�e�z��fd�>����%
�j��A[5��,��=*1�ʒ����=�z�jCo6Mi�LZH��h|l0}�S��n7ўT���
,�\�j���я$�:B6i��D�/��*:��U|گ3f��Z�7�!Z��Me�^����zK�=a�ϼ�';�	g�:	��j��R���Zrs�sφ����[k�O"�\�d���R�����v0�ݳ!!�O~RF�����^uM&g�R��oNOC�D��At&:S��@Ę-|�!��K�y�l��gZ@��ZFJexbՄO>�x)��э���jf�g��H��{�E�;L�U<�qQ�$��̺��k�-� ����Z�j�M��A�si�y֧���/Z��,�"����C�F�����@O�O�BG�G��r-0-�Zgx� *�D����tO�AG����8\y���l���ExY�����v��И���Li�]���)Mdf�:U���F�1ǳ�ݎ�	"�M��9������E{������f����VLP�v@�ÖXߕ�����a��񎘋[\i]TH���Ĉ\�Qu������y��}� ǋ�2K���m�E�A팘E��
Kqbҵ�����x���	����>���9�,�N�b�[m@�h�&)<m���.�{����5���9�t�\0Ch~���/;IR6�Ù<�I8@MOӈ�ױRI�ː�4uf浻s��oD�~�����,��#�$Pr�Ɉ��d��_sO�T�% �-��mC;�Ǵ�����@�C倾�@�H'+�H�X����η������F����(X���Q� �s�Uܕ����Rؗ�l�楺���������	W!��*%H�gjZ��[��)0�l�+~��	�O�F�DUV}��P�+T��F~r^P���A��S-,m�%�fdr,�U���Maj���sH�O�
(3�@[ܽ��D���A3��T��A.w]�������=��o��Q��l��T~4��y�J���L�G���D��-���-�/��'I���m�ǳ�@�2��l�7���67r�l㈟�m�1k������3�?f�HNf��V)бx�O������C�+��X�:�޴��*ňBׄc�%��yf-����XGP����G��lT-7f����iT�a˔=
��mL�-
����ӵ[l��,5ҩ��d�wG���w�3�
��@!�� Fτe�v9T� �,/R��u}���1�X�⶚��I}U�"��]|�m�lv(Ơl��]^���ͽ5��9�N؂�'�M�;#I�f+r�~>�깓��2���}��F`���hU0;c�ʃ��ޠb�|�1D�U�Je�}�/&���1���Y���`_����i�W��b\8��
���:}�|�g��
Af�X�4�fm�,)(�:6Z9r��� UV|6tz� )7��c�L;�����)��iWdIQ+��+յ4J�~x����Y�����%T�&_�T�u�#u�����<0q�y��-�X���\�h��Bc�i��(�FZ/AC�k�BƦ�z���Y&�����g��VX���\�Cm�T,Hדq��]g������s(��AM�����DS:�nAC����=%\ң.��Udj�O�g��ZRُ��	d?�j0C�.Eu�S�vvJx�S�rn�*��d#^�e��	�&Ku�h�����r/��(� =un��+yOw�7�)0U��8E�̈́{���3�I�
�^�x�c4X��0:�K̠��*\߉�'`B.�̰�taG���h��I�0�D:���Q紣�G�J\�@Y2\y:�f�q��d�D�d�ߤD2,�at'���=��)�+w�H��!��<w���w�Ek�RC�j�egL�t��Rote�K:��{��XS���M'��%�ӝ�qy��D�j���{�-��H�~`�hc����.sx����񀁄�oݣB`�Ի9.dW�!���佽��G���'Z��<�@K��J�yȟ8�\C�v@R6�����ʧ�rA9-�=Y�wY�>��6�B�h�/��Y;٘z �ju	\x�$A���kqO	Z��D�Y�+eg0$C�`�ё����&iwa�*���X�sD�0U
c�;B�t<{#3�)��FX�I�/��wR�Y��H��+�S=O#�5[�� ��N���f��a�׊����*!<�^�eM�0Z�"�B��\+�[2���BD��o"�:�*8-�/��aޥ��SA�55R*~�`����G�-���G'!Z_�
clCf��I�aZ��8���Ҕ��?���G�V��>��J���R� ,�j�$�)d"˪��h��X�p/-�r�4�~���D���1��&�H-F����ma%p!�iV$@�h�hR6��jBR�h��=���'ǎD*�*�I$$ΰI��;�M�ͳ[ʴ$A����O�����O��Pl�p��T������$��d���Ͻ�����ܾ�_���M Ģ"��
��� oMשe��qEÒ���B����װN%0�{��D��S�8V�(Wy�x�p�8�˰�t0���}��y��bz��-*�8��#��pO��T��<��D0J��k�B0�H��=}&��viy���p���x�u��5/V�0�욌S�a ���k.�1��J���u�n H��f�t�������d�2}�� 3n7��8ۮ�L��Ƕב=NI�SE�#�[4�_��1>x��n�H�8�
/��R޾���N)�M�����?5g1��e��O�a&
�2����6::F�/���5=.�9�K���B��<��)ۣ�	�A-����I�� $W�AM~ލ�D��t���i�wJ�3H^�)���G�������\�����?-��dx���jN���'���n]Eu�
 �՗��b����P�t���(�w�%苀�z��ᬣz���9|��������'�66P;V�$T�676��f��b�oϧ��S��Q�e!�Ym���f�j��H��HE6?K�>��H�Q�8T��H7ki����:i�t91��{6˼׮�t.�z�?:us�o~Z�	��nֆr$�E1�0,Q�o��V)�����2=~��Ef�х
�Gԇ��U�C�9�c"|҈�ţ��s�-��p� 8�4J�g b}JJ�`�>e�m�W��¿r��i2�q��*X/K�4
Nb��I�E���˔�V��M�K3��֦7d`!2dO�Or����Nv���?O�>~��P��Θܝ�b�{�̞4��9粶�H���K����%[��TM�t��C�֚@�'�;.	
_��lpb'���]A(p!Tͼ�oSD���u��g��fD�Z!&���~1�ö��1��gx����\�l����}��ab�PB��n3��1�����p�FS���S]%�M��K�#A[��/���}PC_b���ڙp�l��D�gI�Fh�=�v3�78�������	[| 8w�����A��]��zg�kU.[�~�r2ѻ�������h�s��4���m�n����K�z���OQ4]{�H"�Gz,�X�����ck8��-ʄ#L[��^�(r
i��� r��j 5�����J�I�t�c|ֺJ��U{��NF,�D��h��� �cBV�F�`C��c�0���}�0?�z�O��`��
Y�g���e��e���E�#���SV��.��w/���&��)��s�����t�| �w&��c�ց�Hչ���V�n���ݷg�������YHW(�&<2���ds4�:�kl������=��5��C�N=�gS�X���v��c�""L��셓%��1l��O{?��lN�v�j�{eu�L�K1�b`0����LW�����\���Y��?BH�;�`_eF���!(-A�l��)E�9��uҜ����j�Х���+�ܯӗ
��H�ɩ5�Q`x<��<n���'|�v�
���J�� �G�f��O!�,� ����L"�)����`zo[>H�A�6����ʦN"Q����_tߢ���(\�h���V��3-9"��q�[