XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[M�t�(��������k��p"=�ݮB��oQ�@��p����#��τ�_�����6���K��@�@g�L�d�%[��!�,`�ê�j��VB�J�%9f:��>��@�?�������gG3��=g������X�{K�cn^�|1r��u���W���R#�4�A�b��@��W�����_��]�=�Y���~�ڜ���|� $�F��X��s?P,�t{!F>�&��A¶�
�L�P{�.�5�.��O�����R���J�����;Jqva�-�H�)��*�<Od`J���
��r��
�$ڛ��7��L�A�',�U(�^�	�Q�x������3z� �=p�䱆�,��Բ��*t��M��xXg���j�c0�%c��L��ӏ_�_D�M˒D��*���1k:�� �����ͣ�<q�%o���k(8�=1��Vx��ծ��W6���5c�F�P_���z)n�{C�K5_�	_k���=��ľ5=)W䔺��`�X�j�b��c�#^��nOv�/i{��n}�{,H��ȡ�a$�d[�IpY����5ԂTY�|��+k����O�>D_R�3��c7�R~V���bm�
�PB0gOI��>��n����
��>Cb/�˔��+PU
u��	Q��C9�a4s[#���L�G�1}��E\�0�,�i�^��(WB����G�
q�p2%zy��}]�t���4_��Wt��1t/������!��Ap,(^�R�|������`���E�m �Z�/�XlxVHYEB    dd8f    2160�]���+��~�,���jƙ,~������K��mC�ŲǨG�]#��X|�+'�W�&���7����6��
�Mހ�"V�w���1g��zw�С�0��/�$`����d��R<,r �U�g�v�iR��RO��y��xMk)l7	n���9:�����I��lx��W����m��Ř]/�.�ؠ���c�q'�/}�[4U�_\�R���מl�t�u�߰W-]�7f�Ҧ�d�W?W>D|�2uٰD���5�um>>�~�;�71&z������ɩ9vR�/?�� MZ-�!��# z��>K��߬�\|�ܪ�$�ᣵ��M?z��y�8W��^p�:����^F���G�)�� >z]���c�5��n)������N��Q�2�� \.��;����"��9
Q���;��7B��"�W�m3����,����������R�G���p����I���OwKp:���nf�6d�J��,�̄x2A[n�����f��n�������R��'�H�= ���1h7B��E�K@��y1�i�djL ���c�e�m�K��jNK��|�:>X�)T��o��߄Sh&�	�Lh�`�q��ǧ��� �����[��;��r��"�����G��n�u>?�9E�I)F �}	�e��$�H�t�i�Z��l@�b��q#�.�k�1�čLsf�@*���4댷W�^��H�<�l�������kؕ4�`���J�zQ��Sk{Q��W^�!(R�R�64J�Z]��������;��3���A�����L���I�'�fm�Ɂf�C��>���tb\eE��h^6��ߝ��p�G=�).'z��6b�g�q��4M��!��֜ݧ��4K:�9 ��P���6L�d�w��o��瘈����!K��}*0�c�*XX3����ċF�j	T�b�z�0��'��a�:A�ӵ':�W��mL,*�c��|&6^t��HıH"z2=���|��}`������{����$�B���q�{u��톊U�'69�ؔhD��2hC��r��ؖX��٦z�N�������ǯ�r7ZEWS���v���ɉL��~��xH2���K"�Q";݌vY遾4��|�F0|!�1��bmìA�"�]J�쮷@ۏ�l�y��&�c�y�%Փ Fd�ԎEI���u}�|e��7��FJ{�a�^�!Y�_!�雺U���_�'E�[ <������.��Ђ9$gC0պ��]#���e%�J@��+4U��0��9��K�� �&��֘��Q�%bh�A�Y)�z]Qⷒ�ҫ��+�G�)?#P�x�j�n@�f�f/čC�ݯ�R�����4�,Y�b)6Ɨ�i��5:06�#�9�B���$�Pf�D����|_Dz5���1yb��	�`����b�e�)	����٘r+X��R��d>T�J�G_?�?��L0]q�{�)�5��`Ck������;��b:x)�f���1���'�T��[���/��̟����d�}����,�f:U��<��S�Ƶ�յ
+��Hn� ��4�L
H����3*U˲���˙��S��tmMA�>"C/#3����HqJa��� �S$�_wr��G�r6�_V�v�@*�z�)B�WL?m�?zǦ)�1n3!٘Osi��?N 8�5�.���8�k�tRUX��C�Q䤟��E�9���/;F� >�6�#!Ŗy�zϹ��Os��N$} U��C*	5��o����F�7�+������k��%+��!Wu����-@|�1��u�?Ê~�[��6�q����+6�c�֥�*��;4�Ced�薞����5Y�Il��>B�Ȓ%lgD���2��o�����c�Q�y�Þ�/F� 
��E��,�W.A�d46Ƽ�@	��Um�8@-�3�5R���f�6loow+>o�� ���I��1D�7<�����-R�2�n�*�t�"�k����pb���Ta�Te+�k��v���_���J���A�mdlu��<�c��&K�+dy��Vh��K�	pd��\�j�з�H�^$?��&d\���*�Q��1n�ܚ?;I���Ť�؋���o/"�����aj>��K8Ԛ�ڐv���ss�^V|�xu>V� �)B�,��`��詣����dF�G������{v�L�D0��x�OgN]�a����k��B߾S �[�Fb�ռ�0N�OJ��M��Ez�ٕMy���)`�E�^0�s䫎��R㙳_��3h|���0)sj�t�'}����h �L�N�~&�dx;H!��R���4�%��	+N{�T>�ְ��11[ϵ�!H�V��x�x�,$/d��i!�b,���z2��ݸgsUDI��	�.8���K�t��=���aюGP҇wY�>s0�C���V�l&eZ��O�|$�N�U(cZa����ʵ���ge"�6�Eb%���÷*Vv�R�dկZ��cZޣZ�ą��eR�i��mz�7����7�s��~Wf�BL]���fI�����Q���'4��; �`=p yg�[v��}�)��R>��5B૽*���=|Y�SL��½a����~L��{��q���I�Ȏ���yē�6�GT���x�\���i4L��l�z3�噘~E�d|�Y�_�	վ�Nu|�9} Ƥ�Of0G<:��������������M&ҽ���4bw/@z���G���"��	��]&�,0�%wC�q�-4����]�f(��V_r�C��!V��J��1�.��r,uϮ{'0ڻ!-uoM���d($m<a�y�c�nW�h�.U[[s��l#\_��Zt�@�!�
�G�xI�mT��$6tN��M�=�OLk	���f�(��UU�����07�F��-G����Ae¼L?�Ԇ&��h[�o����v�
�ww�3�ox��֚�-�� '-{s�⧭^�g�\�G��`��3���C����R;
�N���i���X/���RpֲO�&AݠF����9?cJ�����s���,!�(HOC������9�K{�R�e����GkC$�tj�k��x��*kS۴��j�� �	��U
�ܮj��@ZçB�x���q|U��ͻ��Xw[��/�x*3R;yܽ(ݨaL��U'��Ko$�2+T��&~�8�� g�S������vR�சQ��������	/� �J����+G7�Q��s�zQ��x�����`��5��t��7O^�bS½��W<}�
��d����Ը�(���xt��e�<�[��)�ͷ���c4�O)EgVf��8���W�M�?�S\~�
��n<������#�����g�M���ۊ��k[�j�ġ'��-�Ă��?:e���c�T9��KmT������J���B ab�~�d���Uv�K
.W��/��-z�[�ץ���A��"8�n��W�oq�Q�~F�;$���������$xk�%@�ܪd�� ޯ����Q@0b�Bu r��j��=p���B�&�]�Ta6�`H9=d�]t[#����ؓ��]���1�{�F��P��XI�ǶWk��;e�S8��7N*���B�Wno ��}
N��R��|hb�j�Py(�1m��N
Tj�C`���ٓ�y��ݖ� �l)!I�;�%O���N�<���:P�rt���	�o�M�fAvZI�>b2�3Ի���-dV���6ģ�Q���?'!^H1F���v���Z8h�2�k9��rm��꒬�����hk�~umJ��Yu-�Q���$|߅͖q}'֩)|hjE�gxC�i^�{����%�V�CI�h�	:P���(�:og��Φ>��8l4
�:��|�Q���}sЗ��;��t_�ɐh4�Ԥ<����ش[B���p�o�#���[�9۳\���w��E�o�9�3�4/�CI�URb=z���Հ��]#��?�+Z� ��@%���cE�1��9�[�p��4����/:g��J�ŏ�k��=ٷn����ҍ�
��&/��3�V@M�E�+(0W��M_��"�L6W�/�ZYx�Ot�����6(-�{��I><��_������	l���f J�h�#��+�V�xo�3��M�&]iy9|4����zip%��(���q�pH�s�{���{�M��{��6����~��N��şI�Fo��s^*B
?� ���oN������|I���Wkg�u
F'���_xz+�Z��}MR�d�.8/�)�xˉ�D?��"޲�y^��N%J�"y&׿ec?* L\�#�Ѷ���b`�h�&p�Ü�^>�H`{���ps�s��#2
�ٗ�p�o����U=�u�=25�d>D� �4�gv<�-zF$eD���`|�;��rMx?iw���y��_��C.�rᮖC1w�I>x��׀!#�RY���&\�V����qv_�&%؜����ج���(��K�=�Dߒj���}F1�]q.C�N���}����F6�����a�_^}0E�i?X�X���,g��ud:8�K8y����<N7�vڱ�̴���X��}�����{���g�[��o�=��K�Ə])P�Fb�5�\��H���S�V{DJjP��}L$ Ia�;���q��_�` >��G���;���I:g��j�w�%�20\��WZq^����Z�ѽU2�����7:��d��Z<��$|_�M��4R�@��Oɖ𠝁��-,�ܦ|���9��;�}^����v������8�*g��+5�ߋ+���PV�^� ��>���4yK��60q^
��+�A7[T����2!�����-lZ�Br��e�C���z_�l�(Zt ���R+-N�K��Iʂ����g[N���b�9@L� Q�f��.��kۙ7p~��X���}�+1���%�(ɮ��K`Γ��"s��bpS������͜$/��k���f�ZPDV��*gܹ�+��+�g8�]/N�m�YV�n�ꦒ�+P��-�i�[��JGP�vR۷`�<g�C:2�� ��jnh��K���_=�'!�ף�)ۊ�-B�- �7Ӹ��_)�ғ�4��ɹ�D���Վ�D�K1N��� EaXF�k|klP������7���k�p�^��x��dԷZ�y���~�L�Gt_���E�L)M+�x�ˈ>����%&(#�2�t#UL}�2d��G>�b�e��M�)z�z6�џ�웋F�bt����ȫ��Nz4�5�Τҿ����5,�8��h�`yl�$F���	����<��MV�Z
[廷��!���l�tm���yZ�vpM�}H�-�!��x��ޓ�E��7��!� �vk.�"Y$Z��Xi�n����5�E�kN��C��Ֆ�3ѝ��]G~�.Ϟ�`�g��E�ӡ>��a/���A����*^.U!�0�N��
zer�i�� 	y���O���a�L[o\���u{�|�b�ĸx5����{ 8�DZ8��rK�)X��������"�H�+���������e �;�yYZ��lw����7�Ozq&&�^���v��T����|�͠>��G��)�|�+i��]M(���i�%N��lgo�9�8ےO̳V#�ۅ������牎do*�G���?��pog���Z��.��8��<t�+7�0vl�đ�pe*HqJWND��թ����%�0m���=k2{�"��� �bFz@��Zb��&��t�kg簉�8u�A<�?���Kl@:~��5�F=��w���mڭS.��L��>�g_8t=>�U�"��3kvg�>�8Ē2	���b�x���P}Iف��؈u�J�܅ϭDm��^��#����J7�;���b��	���(a��RԄ�>��O;��=O{�eW�OE��S�%�, �����D�7�� H�,�PH���m��R'R�&�ϊ�~󆔣���7�YP�ѻ���^�좿�Uy�A��J��.��h>��2 �ӳ�i%��� ���U����&b�V��)�d:�g?HY����!Wm�����2�r���
[�L��r�e��뽅5�Dò��M7\,���K��;S(K�w�v��5��5R�s%jl(ã��AJe'~��T�UE�qKU�>h/�ޖ��|U?����fT/Y���S}�Ћ��,�np��^%�h�}������b���Bb7�.����+Hr�Q:��Y2O�7��ꢽ�-D=�>:pzYh��(M��� /��a�s����R>�Z���OL�W�V��rPCx�����$��߃��� 6f=��% u�b����BF���Y������t�wR�)vd�\g�g_�bU8=���$MjǾ��7-	�fF	�����ł+	,���&��#���6z�ne��z)H�"O��)%� �˴�W���M���Đ�����Y�����I�~*�F�a��׶i0(��:skp/92� 6B�F�$�Nyi�{A .�.�3�35�-���S�!#(��n��� ��*&���8��y�H�qr�(D5�����O�:�P yW�'<��UaM �.���l�h[�m�c������e2��V|,�w����v������RC<OEn��:��^�^��.�R���~�>sÿP０6 ˈWO=w�R�tm�k�Q[u1��hH���`����@Dj˼��d�U=�7sag��-������+gW	Q�b]Go��~�N��]�;f� 8�0����u�LD{ Blԙ���@ٙ���L��-bA�V�6MYmj�Kb��ᡲ������~�޶���~�����G/��Ti]�����~�%kK�,�'�~%�=f���D>�ĉ���Mfx���_��|�#U�X����xIB�iX�V�3���g_o�����+����o��f;M콐O��.Ю�C�� � >�:2���7��U2����2���{��懦K�sI�hw���� "4xqX��9վ+6���rx�ކ�9����!�9v�7�sM��������^��w��hx��C���;�V ��?��W�t얂[FN���vaMԻqR5w��Eŭ3%,s�a�g�~���"���YMYV�q�5�>"+˖��KB���	h7�5o�v5#��*�Y�s�#0C���.�i�)}�;�2��7i>�ߺ��F�|v^T&ԀV��q��f���qQK�CG�/��Z��218��י�]�Z8{��ҥ	��t��y2���\l!�
���$� �Lr�>����߶}��y�A3O�s.6�қ�Ӷ�v��8�W�/oi�P�����~�ސ��*΁l��ݘ)�Eg+48�z�C�q�Bmc
�z�hE������@���a��;�H�Sj��:� �����E���!�@�Vǯ�;��~��7��pV�0ZOz���q���=�4&�0����������	̢���*d?+6FV��QS���U�� ��ɱ�b�A0�Sxߩħl��L��_�zլ�)�'��̆�x��4V���iDW2���oFӻO:�,���f+��D��w���R���&sع F%M�uW��.a�9�-�VON40���
���{�2JZ�v
X��������9�W�bsC��7f���.���5��i��z���G��6�]?$A|��+T��z��-�̤����r-7�<!`/B A%�,s��XG�IR�|VdMi����)\���@�#�锂�ث���tN��Q���������gXD����&�Ӧ$�kx���?��N'Tj���~�Ǜ����A*l� ��9�j�r�.*kz�U����YC��:�͞���dc� 7/�^�Δ�U���[�����B۲+f�T�]W_:�b������ˮ��!����)�� ��^����(�M�e@%�y1��s�qiȴ��-�}sK˥�L�s�~�AO.��'?���._��ڇ�Y/���0&��_�{G@A����� LT���S��p��(���j񫢿��8н���tH��Y\������s,rҥ`�{�G_j�2����J�������J��L�y-I�q=6��YN^��E�n��t;���1��U3��-�+�r`l�'(.��,�.��&�_�b�,�
P�杠y<���hj�N������U(�X����s\{?�
J��BMS��UzZ��ѕ<0�>�"U�j�!k"�imH�UA�����;2�Y�}���?n
����E~h�����(��������[���1#�6�-bp�/�nct�x8N%#l�
��HV���XK��D�zb�F�ݔz�W�cix�f�13��?�9�^�� [DI�h��Z+_1���90��Hk�!F�gYU�܊w̤@�q�JRM���l�.���R�ul�@'����7j���TʇAj��74�K��x����Զy����0�H�uw�7bzj��Y��p��l�Z4f�