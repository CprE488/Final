XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#��zE�я�c�;?Xi��=o0%���}���(�D�iF�Դ���'p��mN�	���ѡ��@~x.�ʠ�k���!,XN֪ A��9��R6��o�FAn�G�wɐ�k��mözD��b�z��O�#u�)ow��������h�a\�$��Dj(2�L����ռ�J���2�S5eD�P�������3H�al���b1L'm���tI���QR���v��۽0!+"��fk�4�+]���-�3$V�Rs��A6��薠rF�K<fh�w��G�L^6���{���|��~n�N��Z�;�ѐ�E��I+"z�PW���5������G+�Ć�"�����)�t���D�������ǀ��ŸF��+��&��a%��m[��Af;�Oxv7��9~]Fix�:�!J%�B������#���*f��aJn����H���$sI�M�;3-�W>��{���U��9�p��ZN1#z>���/���v=�:W���W6��_<�	+( �s��E�Nu(�g�������ZMp�ԃ�۝�U��0{V{E��r�;��Y���X.NE�z�A�[�}�	�Y���9��wt��V̄��b~M.iX?�W4e����-G�d�18�}�Ĝ��(7�5␿״K͕:�E͈�?`)��<�l\�)9g�yT�>ed�f׮��\�dOb����Ȥ�q8�o�ݤ�u�ȠpȖ����p�\���GOe$@XlxVHYEB    b3c6    25b0���A_�gr�(��W���Z�#�0 az��N��������0����8pB��\����F�0UO�]�����e^�Rڎ�s�1����V_ ����{�����u0#g���9c��ssP1�}�m��(;KT�d\��3�TX����_J$+nuӣ�\��!��Qi7e���a������\�OCh�R �(-�1�9Y��r�Ȩ����X@`?U��� ��c|5d���[H����1�:��zU�xt~�Q�UM���hX�B=�HP�?���i�w��LWw�)uV� y��UH�>"$9H���S����	�w_dy�{���6}+�������Ű%R}0w'�B��16��;Qm�#�\~��f���p���]�5]ؕSI��Ԉ kJI�[Q�_�����6�i��9�C{,|�2�b�Z'���#V�Xpo��?�C��	��Ȕ��[�#<���5���U{���"�u>f���}_>.e`H�|��T�n1=�Z>��ڪ��!���f uqC�2����F��F�%���B1�}#��C��&�����;g��@������[̩YV��O��,�)��'�7� g�����)��?*��㰓�*f�w5����ᕗ�C��7�A6>?�:m��hd��V�̸��Liõ�5�vJ;B>�G9VP �V;9Mu�.+�����ԧ�E4.��FWއ���{!�7O6���* 7,d�hFI�?R�Α�\���G��O_��P#A���&L�5�y.�=�t��{�tBSg���Yf4����Y�ѩAs�I�&5Qxvaϟdn 4��/C}�Q��C�'��	��~�Z%e9�t����g���)��l���O�bw�5���j��3u��H8�Qq6�O
��S��|E8�#��vJ�i��
�B�T��E�i�`~pw�f�#���'�����#D6��$�<�2ܻmQ�?b%YtS�?pD#P�8	��C%�R�5&�X4�k�&m�ǘ�.�7i�@�S�Ns�����UֽYwF~����64��'w�����!�AYU=�Fh(�ǅ;PFGB�6`5�^�ֳ�ݿO��+.�b��`!>	��tǡr��AT��"}�F�#�yzL,�]17��P7f������V�IAӡ�#�K�Q��E9��I�&^qQ&��x7}J7���(}�Oƹ�(���@�7=�Ԩ���-��EV���O@�f�V:�@��6��;o/��ʓ�5]E�St���� j��@fY���UBHU,(2M ��|�T%��y?M���8��h�6-'b���N|DM��юߘo-����3{�^�5��d�f�!H#�
>��bx�&[�_�L}�I`׾�'��ä����~����͇����(�����)�Έ���
�2:�TE5�g�������6$�u�e���ʒ��N�3�y������{#�b]1*������AH�Xr�T�'�4��䟖y�X,<۷R�߽s�<�'�+S��NBI�6�K��[�FU�N"G��س/��x��ܑQ�Q��Z7�e��o���8/�A��w��6^�#V�̗����]_��V8��F&#>�˽ي��z8���b��o�yb��%�$tK�U��d0H�%�I|�J�}��O���ɬ�*r�ao3���۹��=^��%�^��me�E)Q�+uHcu�0��L�ר�6�֬m��-X;o��	�m��K��f�
q9cSBL�%9����I��G�����fY��#����gTץ7�Re�R�݉]��H`?d�p��\�ٵ�dq�{���gunu�"��ȇ��_o��bǽ�+,��i}.�7Fڬ��
:m�<Y�|�Ÿ8l��L+;�nB�\�YRQ=⩑8������jS������+�A�$M�t���>��W��S)Cw�C�Q�ȫ\
������|p����9�U���e���+�D������%�T.�aY�`��t*��ą
�$(���&�d6����bF������#��~I��� ��!L�`z�y�?�L��Л���K��`Q���0�ɧ�+�u�G�I�����n��Gv��� αF1d����L��b�~�<y�8�\����k �?A�xq�,��Y�7W?�+���8%Me��>E�f#����e����۶�YQ����9UQ$bi�q�A^ZM��f6��Sp����e J�	G���'�y������'.�Vo<f�#�_�'C�c9%��3���Z�a�@��g��~��X��@#!���,��jK��� ��U��'��H�e!p-��� Ӟv�0<�Z�?k�#��`�.��YWCl�7V��rP5m���4"C�萯�q"U���<�5�K�!���l����PQ��h�&g%����ygy'�����A!c��#�N��M�OK0�]��}l�
�b��4��.�X�K)ƹ�͑/�@Ѱ6Դ�)0�8--���<;���b����� o�n��vn�I2"��l#�6O[�x�u�&I/����}3�zwå�דg�Z;s1���u_�kcG�r ٍ�*�~a��%V�s3֨g�c�i�3�۫�h�
�$�Kူ��̑�c�O/4>�@(��t��hԾŏ��,H��}@��O�������Q�(O�J�Z3a�R�hu��I]ky�9?���@��Zz�>��ǳ�*���VHaXl>�x��x��k��f5R� ^���q�ř�=t���yR�ע?�Z�����Y���ӿ��[G69a��pk�4���Ql�M����ϻ�*G��M�r�Gv��<!SfX����A��-����t�A���BYW�2a��5�]Z2o6���'V�˴�{���O�S�ۚ��'��;*�h�B����]��R��	��s1$�\�Ly��r2Q��HA�e�X�#c����;g���nlχ�ky_)�J�v��<l�<DA�σ�`�j\�^;���ڲ����Ud�dE�c�<��oم�E<���WL��)~��{�5��ƭq�"��p�(� �{:����X4�����o�+~e92*���GGX��O�
�h�Z��֡f�X�>%��?�e��}	Ǟ��'+�9&��\��ŪG.*�4���7�DQa�:B�����KG���J'�n�ٶ��f=�?b��� x���Fyor{����?l�f'3|�<�G�$_�Wf���VVM�q~&� R�w��Zsq�PbW��39�����]K�P!h#�y�\!W��bj�Ċ��� /��#���y���+��*:�f�J $�9'nn���>����ʎi:=!:����d0����{�>1&A���vf�:������ǖ!��b�3��[O�y� "L0��s�T���~ԥ��<I�'Ne926�S
l��TA/
qLߚ��wt����Ϻ-~�ž���@r��e�E��3͊ �fq��П���_���{����w�n 1��w��4�OK����yG�9J�u�[��!���O��Q^���G��*����Da�)��&�T���=,�!�y���';�z��i�fN��_5_-!�F���N*=P�J�y����ĸPsJK��SHK�d���2|�+���Y�U���E��Z�36
��|��b_��r۞D,���v�,j�a�;���Aj�`4ĳ��XWNG�g�ZӆpZN���
�)[����,_�@a��B����#-�-ϙnY�����vzRmJy�tϼ� �
�G#a�xL���T¡��ft��O�z��m��'<yZ]��?_ѽ6LѤ�;��%XLV1����&��X�n�Qu��E�5\�����ք#��O_��(�||v��<y��?m�Ie	���ϼ��ޛ~�J����;dL�	�����o�:x_�1�8g�<��)m$��C��F0|�T�0��V܉���4���h٫��n�BƳ�y�qn@?e��R�k��.vD�X�6�N��{wk�9!�m�%�Of�9�� ��Dܵ[�?�����-*�,b��,%Y���W��/�Z����r��/W�MC��=��;ǿp]�}`�����B�Ƭ����/���#F����t�����8^\�Y��:G85�o��m#}��Ka{�;���3��16��r�nޢ�s�rά�[(��\2�]���|_&ۄys�����v�������%�G�0��bp�TU��k���Q ��fcf���%"I`���
���u�
�2.}!I}F���mo �3s��I�A��W��1����f��H$���Y��!*Zj��C�)���髤)�����������U�WOE`H�NA�)��#m��i���潄 ��?�����b�W��_<�\�w�L�%� %q̴L�w�T�{���h�"���+6�)��.���Ef���eV9���w��}�7�f仠��t�I8J~�ӊ���A:�r���U_0J�F�|%%�j�ʲ؆�JGŏ�p.��z��HaB��"�*a�����}ΥS����Q�7Gxmb��ׅF�i�9|�
����c|�Ϣ�r�"e?�e<�Ɋh)����S�\����jɈul�����`���%M�%k�P��F�~뭤�j��+��	�l]���PCt�bR�;sm��$Ĭ�e��R�Fú�?C�T��wr��ښmOk~�H�����WU������hCvm�ר���j��:j���Mʫ�h��嶛A�;�7Ğ�4!�z��1���x�����gd�%�Wp�����U�v������?K�;.ƛ&�Q`�S�H�r�<�-J�Cj`���p�>6X�c!�Wiz���S�GZ��ws�;�Ѻ��LIu|������
����˫���IB�M���wq�\�!�JNr�蜅Ť[��X���eܲ=�?J ��h+t�~ӳ�>gc=X`JFZ\�p����S�7���XE�U}�JҦ���Ո��:/=@l�� ��UM|�Vv�(����-u�I�����mDsA�ǔcI�p�`l�~/�(nox� ��Z���U��FG.w1Z���J5#�_if�;����t���s�m$m��nw�7 ���-�	?<3OL�/�Q���}9H�q�b�Ɗ
�7�O�)��!���)fȖt�D�6Dh� CB�Aj���Pep��pL�b�~|Lx<��҅����9F�}��u�f!rI�KD�q�}�ھf���%�����(7�Tw<���g��>��m��˴������͞v�@Ңu]���rgklp.�h�I~N�>7ɂ��8/����/+fh�����d,;���q����Kc.��*�XO-��̸i�3f���&4��?��O�]���	r� ���{�����2���b��B� �K��Y�(ݾ]f�[��h^yN[J�8���Gr��v�Z?���դ���w��5�_\��IRJ`�h�B�ر�b ߃�; �O��[������*����v��3�5����6��?�f�9Jg|l��tGW��c��{1i�nR\R����Vn���he��:���ڒ,f,o�r7y	���UI�ʳ3�a�g��E�b2��O���)�� �����q~��R��S/	\��v�Y������5����$v�S �/i5�!�N��o64��o�W<J\���Ӓ�f���,v�j���lF�^p�G�� �Ssqb���ɋV)��0Q�0GyG��k�V����I��:(4��h���Q!Eo���Q
͙+I��9]���]�n�}��MF->D�#U�Ǆ��B�>�K�{���ZT���߸�;�?��`�c��H� �r��bw-q��%\wUF��4EJ($`���W~4;ǰ�$m8_T[��/�/zgGF{!���<U^�	�U�U��% E.�F�>aR򭮲��\2g�9���+�{/�ТC�o���䬜��^oB����P����::=l�;OZO������R`��Y��e�Q;1|^->s��F
��W/�*�Oc�-~��ϗa��r<=.��;#�ϟ�L[���� ��?�ʁk�U}�eЍ��y+���ۣ}�� =6�˴��)v����7�h����mP�OS�Rxx2���R��a����W���z/�&�U���[hB��ͭ�A1=�4�d�,�o�"6�<Ⱥ����ROVKB�?�����_��c&��WZF��D3/и}��s����5�?;�,�D�9����%�+X�3po�Xi]���l�bqe����rt���N$�n.f�۝�Y�F�� �ю���c�A���~1\y�AqH���M��_x�~�F�rZ6�G�-!<qNA�Ϛ��T��pb9���F����&B>d�MC��f���1Xm���ܗܵ���vS�U��9���~�����n�̨s�i��R�a7���(��]J�n�dD�Z |sM�jP@E�� ]��!�����;�lwi��x�IHC����)�Bm��K3�-PI��C�[E����a~�%��ԛR!Д?@�HU��FO��ć�f�-.����k���Ϭ��)�}��� 
"��������`�O�b��e��X���v��.s�(��.�y9z���#3�Ď��3{6;�V� L���'|��E�m�������q�6 
�y=��x���%�r�w�\-�@>�|����$~(s
�))!���t�j�@Fѕ��H��3�|?T-����zb�n����J6ݒ�a�;������Y�tJ�RB��odI���`|�R�GW5	��L;kW[H��ˣVC�.c��.���uw�EdD�O�:�yPҋ�x���E��l3Z������+������n��!2N,��)֤3�a�t�e�����y���SԬ��'|�֦xsx��s,r@��n)�)}>�[ɀ�ǟ��S��Z���R]���D�l��j�Ɂ[Ie��S�V��#���	�@��������˃_��oɖ��o�"/bI����U'灜1|%|x�3����9(��F��we���|U����ΈX�}p6
h�K��`��6�z� I	���萒�3N���a*ry&��־�q���+�d)�U_��P)B*P)�/������e)�7�KYHQ����8e52}Ю[��BR���|�M�X�Hwr�6��v� Z�q�	�v�ɉ�G[~��+���)b����x�Ԑ70� `��i$ѫ?<��ٷ4Z����	��/;���TP۝^[���[�e�4����ư��΋�䭑�� c��]�k��l8����o����äg���S\��:��FfN�������b�`2I��S�9C��,�	�ݵ�2��%:�L^�*N���9V�A���Ki��M��DWA��}YꥋN
��;�>0���?�h8����>�jSۀ{E�9��Zc�dR"�v�֥�d.��.�h�%q5�����tE�9��Y�,lm���ڥ��'�]�6c�z�Qۅ�J$7�3�?͎�x�+Wp�Ta�*�1[�8#}6��ot����|j�u�d�(��$��w_�tqJ/ŵTV�[-�Yih�&C�ޑ�u-f��3M�rN�k����s?��_T7�KMl�G$}DG�d�[�}��].������<f�ݏ^�?��[!�9}���dbVk�<��=RQ?9�� ��L;�Y_����Xm�q��N�/�O��v�g[k.O���]gS���	3$b���c��B�����uoO��2l���;�`J��8�ݨ���RJlR�B7H�m}���чbl��8`�ܱ�<imEk&Yh,K��ԓa���Y��ۍ0�S&��a�zC��`ƥ₈N6�<�9*��,����&:M����{�,�Sj�JL���!�g���v)�H�d��骦+k��w�IM5�◐p$���HG�����B�\�3�^��_1+�থ���fʺpnJ��`�'GkK���E��~Ȫ��5kR��ϧ}�C`-�0��Kd�#[��}<����'�����/0��+n�T�l���yw����q���
nb�lx�}���Of]�� 5�l$�",̦_�TT�~���!�i�v�U~$V� W��и�i�Z�������`��)��x��*w�TX����%|n�J00�����yc��Gkreq"������XRf��ƴ�;�G1�dY@��FSKc,�y�Y�OW��Y�4|��~�H)_�-� ��ya���9F��*4z&h�n���rx�o������VL��H�F;���9.��'GG���v	Ɣv���A��n���J��^��/��I�CJ�=VP�#�%�J�Z��t�����+����lfĦl^��h��9���}����
���E���I1��&	�1t��p�\{�U���:��Ib���2�R�Pڌ�ߥ�S�i�+��l�uA�=D�q�$҂w�02/͸Z��] ��|Du�k������L�q��VLM	ԧZ��:���^D�w�3|�
�du� j��e}���N��P�`3�V`���ܓ�H�`¤�?�a\�/km�ߎX��b�dy��d3�ul�[�0�)�aFd�h�5�3���n5�F��}?֢��3v�V9LaȪ����}$���l)�!��SV
�tB��}!��ZC^#]Pl~�BU���M�EǏ��3&�^K����nL�x�D���{��:�>�K�(���hgun��%��@p�e�
W��3(u�%�3���ъC��jv��n�ڪre��U�kY�������9&B~Ԍ�/�{�3��i_}�6����YgL_j�1� �,Rr�]䧡�^F�n�*�����oL(~%u���c|��׊���!H���@��9>5��ϳ�� ��Nk��#�M^�@8t�:��*�%A�hǀ4�����#!���]�z��X �}=G_w��;���җ���O�J3ݴ#��oK(%����<#�,�1+� ��{��q�{䠹X<��$��SW�!�i�$�H�*3�8a���eH����8���H�s�B�&��d2���d��h�^@S��7�Y��)�.$d�k����L�G���t�3Xy4j�7=�Ԋ�v�1�ۗ� %j�-��:�=C������)!���k?f�N��A��I�z��$�&y�֊��(�° ��!s�C4���{m�;�9=p4fcۂ5Բn��
��E#�l���o�����b�pr.������t�K��Ǚ����g�rK�X%��Q4�4�Tq��w�x�����]܃o�C�A��U���~�|��jO��(6ڋ-F�gI:0DV�W F�v��w�*U�Kl2�w��1��*!Z�~�?��D�j㮧���i7��U��?���4��P��a�6���%S�F/*�^��^q�׋�x�Ϩ�U�.�D���qh�����+��,���wԴ�.gku��Zjn�����*��J�WSҰ��+�zDc�
��uE��Aם�xu��R)p�iBs*n.{�3�ݭ�ٍN��)GRN,�ąs���r�@~��"H�m/T����U1�5����