XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����M�X��bo���X�U�s�θb"(��G\�9jY.������c�{v�8�f7������s�-M�����-���Oi�.���,�	���_&���f�R!��N7�[%?����,.�"���_)$��e`ZԑG�����=N T����0���"�'	yUC�zB�ՠ=���������n��,� k΢���5�&�k�8j���c����`�n'�M�A5_J;ĿH�u�&QA�o�QRr�x;'����&�����Z�J����1غ0Ŧ����&��-ܰ~�%y�s�@5f*�s>`8��`�����J�f\G	�`��P=���$��Р�vfaԢ4�?��P���:�(�#ŵOXk2��T��f���Yἐʄn�i��;���]�6ܻ½�ZꙌȣ_�'�b�q´&D�^�U^Z��i�� Ԣ�f�fL{+h��#;�R���49��s���_�E8aٗ�^���o����<C�w�/uċ�̰e8�_�:m�b���Z��w]���|���I��s\�pc��Sn0�Gfi�a|��&o�e({���z�T���-�h�#��mv�+�b,$�s��]yy�,OB��"��������)ǕG?�mBE�n�ǃ�ݏ����a��2�|�ܓ��3U�h(U�9�<w�z�Κ�i��S��"��Lz2��-*B8�n�6q�rv�VLz%���O�&�C��~��7A�G�c��P핡�,U�����)���0�e��̐��XlxVHYEB    1853     810Ʉ�f缫��+U��+[��-��2{Gb^W;�]'��KI.�Κ�H��`�:�G�.��3�)������\����Vyq-����!pq?��\������d�e:�(G'Br��(kN��~ �tj���j���6%�9�~th�2ށǥI��뙥��
�&�/����5 �-�H��ɦ���&��Z���S�����>�OzVd�����N��p����]����t<��_�3���ic�}Q����ﯥ�W� +����(�����
D�[�QRqL܌BH+��1��ȿ�ҋ�b�%ƨQ!�m�}	����k�N�)	u���v�F��?x��}���-��v%}k�=�خ�C0K��s]�BID�g�90�f�}���[e�ġ�����w�#u-�G��z�v��ĹrCi��tGV�C����4�*G�o�F���W��O�5�%�^�~�H���sS\�>;�����]�P]���T��z�8[�<��^���@������zC����vD���Á�~��S1�e��]ߘ9����^���B�v[�ԹѾ�>��|nI ��J�	��p�]&B%��cw����1��r�z�ndV�x����6$��V7���z�+��K�[�wӲ�a¤�a'��O����O`�,K�L����E�О����8�5���@��st����84 ǃ�\�q��ٞ����^�ژ����;Kq��S��?}�}�,ӣ��$��=�B@�Z�P^Hh�PI�]!?���,�dq�R�����\G���1f(��U]k/`<"����I"�����d�s޽�g�8�̆���)�~�~�vm�cvo�S�4��j���7;[�ң�O�s6
&��p(c����o(BK�o �-^�� ���yk���~����C�������zS��O!�'Q�O��}=
���X���+"	0: �{�Q�
��:<�6��/Xce-�
sf���+�M<�$Jp~z��cA4Kc�~Zq�kWج�zYA+��U�%�N�*�P�v��C뒣.+��{�#��{�[B�*]{�O$�`��w%k���!4�o���׭{Q%7�+�� ���g>6DY�~.pam�If׽�� =Ā6��?�C�0=�n��NV��`���)��s��cj	qKr7�P�|�Z�M|_W�Փ� #���^ހ��b˒Ƿ������Xz�=~,}�(��%�a�r�Hw�nϝ�/��w G14��j㒀3�>��|�Ax�[��AC&PT��z\�q�$P>�@�PH���ß:�#C~tݣ�!!�M�+a���;`(<?�0Z�+Ī��$k/��Wp���7������+&�Ɠ�:�N��q��8�-ݣ�	�9b\����#n2Ҽ$$*������Ă1�ϡo��]��~z/�
_w�?&z�zw��h*_��+_�(dV����'C��/�9�Úb�H1 ���e�sr	�8�x����u�;��ƻ�����1hQ/�[�eXm�P��@r3ddXBD�����s�{pwS�G*����~�q�U�>�(q�׼A��V�B���h��q��&�%`���D2�u�\����~�|�)�@���4��O��j��X����8���:W���T�1�����xx�H�Z��6�V!Xؽٙ�N��4e ���7����+����?�K���RK��#�O<J˔����W�ec�0ȩ؜[?�z�<�W\F>Tg.}W�xwBi��9��ZP�	P)!R��B�9�(w��E�|f�Ǚ��~4���l'��\:KM���$<��d<�Ky�E^sm�t�^S�Z�sg�&�������<����^��g}(��+1`�E��k ��Oy7�O�f�Z�����T![�}�L�*4G[%�sI��m�Y^^/��P��2k���]�D�`Í�u%H�rs����=fhI�<i��l�����I��-Đ#s����n��4�m�#���h������q�B���a+�k#@�'bB��v|��N�)s��b&��;Vx�2 �(eG@;�O�����: