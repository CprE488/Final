XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���a�/R"�~�E�>����ɓ�/K�|wD��O���[����=�����K����N'��$��52�`'��ߧql�=�S��@=�N�3-9@j?���S���	O�����b�8��pEC�@���3I�)y��͵,&N鬐"�Q%9�IZH��z�}V��=���]�YXTy����K'���J0Vss�/�|b]�+}�[�XC����v`��{~�vwY��P[k���e�NIN�؅-�u�0���n��P��+`�Ȝ6�Ekc���i�������Zo諅�P��O��4h�!P�3��� �l�ҹ�x[~3"�����BDW�xWÄ�`�R�dW���L�C���d�='.C��1��SQx�'��|3�KL�Ԁ39֗coC�Vv��tvl�1�j#��a�Z�{_�:lQ�,M�7�]@�+�$� �˺�� *����V��weW6�Q�x�0�P�u%��LV��_Ƴ ��hh&v�Ko�\e/)،yhw�h�E�9��:��/Db����i��� �[���AW��!�|Q�^/Q��qsk<�؄x�+�����=p���o䔂����kM��0נ����l��iF�k���HM�i�i�77�N�c��:�������܇B֛����8��MsJ��&�Hw��#��ٷ�γ��{���R��^��K��Ǜ1R����.�K���a���D��g6�����C�.ɘח?)���&ɉ��<ͫ	FeAM�=����S��ͧ�F�XlxVHYEB    6346    1790;L�������w�F�x`v�í[l��eM�U-�xcM�Ό-��|f�}�������h������@<S5�\l,��4�����˶z��Ȍd��r�
�8�n��#տL�����MR��s��ۦ?^ ��8H+�L�g�R7� ��G˺o3�@�3����ĩ��/u_qM+��_�,��4IB��}m���GH�Ee�8�=ėG��	<ׇ0�3�r����^���FN��'�d�r̿^�����r-��Rz���r�QEܙd���i����x�֛^�k P[����C��Mr��"�ح�O<�sV�;@�b��gq���7��Z�۱0�q|���V�n�?��)/~͇p��urN[�- �zz$�7�����l����iHv�7f)��=��-�����˕�ů�TF���I.+�x��y���h��WO��[�j�ЈZ-�t���i�|�J6q;6�� ���f�}�EP�OU2�0�X�a����P�{���V^�
�@�:��
�8���W[AG6��c֛�]_��.Xf6���&��;�u�;mnHwu���@�\S��ݬ�>��%$��4Փ�J�!����0�{Y����֕@-@��(�p��o�-�T^l&:�*W`�ɓ��E��0�g�o'�\�o��Y
�~�s	}	a�F���{�����2N���2��`�t۸N0�aY���$#B&�}��R뷳#q�%7O��y�+�~��	���̪-�\�z'ž{H���r���x;_c��p���5�����˲0�}�J�;/'�lz�I��9�W#����h f^lM��$[�̞횭�^C�K����)�D�98�a������������m��AE��p
QTK;��Ս ����C0vp��c�)>�8��AM�P[�* SM��j�Xq�٫cR=��א5�!��� �C�5���I��Ҿ�@�e`>'#�ߐ��5��焪�W��)�g�����k��� 9�E�M5Y�Q��Yp=��n~I�c�:�qj�UZ���͙w��C�7�Ա��[D �Lǃ�g��IK�q�[`v�A:*��Ӟ`[K|*-D"�6��R�����6���9 ̤��Y� H�o��Ǯ�C���֫��W����OG
�Y`c���:�OB��@�E��~~���&(�G�3¥|;ό�h/�D��)����j]��X\�n�� pC����������'|��au��A5oMh��သ���A����¥�X�R4��m�����$9� �d)Z�#�+P�x
db*F��#x�&L"�i�@�	El�����0u�y0ve���4=y�	���ڏ�| ��uZ�svF`W�w�^�YYK��4J���I��i���dA�i�Lu��z�tt"|�#�`����&3��Ҩ��N�;6u&4"��s~��.��{%�v���B�C~��z��|�T���qזz�d8��|`��rD�qݵ�A���)|]x%A /��wm�p�^�E��T���#�'W_��Ջ�;�7�d���8u��^���rU��T/�,�?�c�N��ʶh11#�K](A��2��F��z�6lb�w^	Y���~x��e�~�Gs]q# 92$�aR�*~ϸb���������p�g� ����L��1��'�2>�X��ʔ�0	ݑ#��Q��}�LY$�-�51� >Ŷ�iP�e��YM{��Ԃ�&�8�t&��m|����Vl;}֖`��Fϰ��`Ͽ7-i� T���!��j��5����Q������Ǻ�ؠ�.߁Cy���Y���k�HAV�1d�Õ��a�Ƀ+<V�=D�}z�!ȕ�����_��O=]�99gjU�?�8j���E�q$ek�O�k~�#�&�ƙ:R����O8���'D�i�[�0~�����B�^b�6�w����, DJ���MW���0�G�Q�V�k�f�z��X���m�U�&[��Z�P|���\�A�Ð�G�aF; ���� ��f�� ��KpV��LSf��#���[����)��0G�\�U�$$@F�EC�[zI�%E����u^�U��`"<��u�D�^��!#�g�I��?^��;K���MG^ܙD��e(�P���3�wW�Q�	V`�vǔܚv��.-;�G�N�Kڌ�9��e3^j\��(��8�C�{�?n#�%&�N��;�ۨͪ�a�SO- 4���!��ʐ�e��%�,�K`Mx�&?zZF�q��c���Uv�/�������)�Z�G��/b���ؒ���je�:�|�ۑ�;��f���[/����ޭ���:��������A8�z�S<
9�����I�@�r���Jd�U�5Ǡ߼V�b�������{)o�Z��54QL$%�>wTǱP���Lfk8x-�#��B1�崠V�?��?�Π��I�s�w����r1��>1��cF]���6�|~j�n���.���r�����7�Yˡ��B֐g�MF����ǟ�4'�:�"5�C�y@�)oq�O��	�$��b�黥ѝQ���lpO��&���%���*��gF��S(/U?::�'Q`���x���Y,�"��P)���3�����/鎾���4�����2j��.)�M����Ɍ�C���ʌ9�;�U��.���t�O�����U���u�n�S=	��s��<�
�7<��;Iw�mMFv��g����b�T 0�N����X��� L�\�pl$2�H	Èy'q�=����)�q��jx�Q��N�O�ө���×�NJ�b��{��Ǉ�{�LC-�X���&�;B��������K �ir/���z~o0����Se+AD9��B�ٶe�;h�\�|�;���cZgi!y�����r���x�U�Ec��`���z:46��[��>������3*s��΍��x.�IU@���~�U����o��ǖ���IYrs��	B�\E���'~h�l��e&+nL��{�g^�^�U�����Otl`���xYJZ��I����WN0������lԤpǹ51�4l�*��آ�+�����m� �M�����Hr��GRy'��WRl],����M�%�.!���>����l�Q���&�A��}��*N��	0p��,�0������9��~yM1�x�V�,f�7s�G���&�A-��z|���`n՝?h.�x�?+(��M`R:��"�zNq���~j�yJ1�q�0\�����)u��#�V�7����<����x�P�� �%��B�%�nX��N��tp�L��U�T�g����������� ��˾@=��;8�9��&�Ë��u�*���@34�w#E�s�Zg��MJl�o����G��(c,�b����"��Mq(
�w�t'��"��.���X>���C�����:n:�[�c�/��KɔкH�cb�Kmh���^S��O&�?��G����r�L�o��]�Q]^(?���$PS	��$YS^����-I\��n\K�z<�ݺ�u3�OjtS���|Yʺp�P��i_-\���9S�� �k�&��æs����a�8	L��5���n��>ښ��T�V��Dt�]�S�[�;�q
?����6`�o,��
�:�n4ޤ��q��T�)���Tn�<����AƱ�g�Emk}��Y&n�u0'�����յ@#�����L��܋��nH�[���aUȪ������E�^hC���\�B��ysϕ��?���>Ҋh�P�?�}F�j�_Gh�N?�e�tB+@m*r�|�[L��:��$Hnl�}��*"^���yΐ�98����3f�G��M����R�·���sM��kJ�=/���7��9�H�?��@k�Q���>ڂ�D )��Z�R�(�ٚҧ����G,Z9�vy��Q�g�[0oN G����B
�*UX�$4��ݣ0!�98~��ĠԬ����M�e� sp	��H ��I�Ip�`�x��+2ON߃S$�̎�y��}2�?��T�YL�q}���e�*����@���X���Ó��@�Zt[�؟*�`r1�����vq��sо� �~���-��͌z��"$���;O��'�n/e�N�@�9��-9��wD���u9�3iEp�˒�	����%т��3~[�
�+�N�=)[�KE����]��l3+M��'U5y��|�C�n��X��3��N>�;L�	�'p�})B��H�B*@�P��L�9�R'���5!1��Ia˃�Bm����9��uV*r./��^�?.�����:�3
�Rc�	ZE�%<���:a�s�٨��*
����ˌv� j.�V���V�W�У���&�$`$52Dw�Q�1kcN�Z���3�#�#��i�B�p�a�O�F�]\fl���C8�Lq���t�Г��#��|�^5>Ǜ����V��g�v*#�?���oaR�9!�-�1���/�����8�2�g��xD�m߁,�o��3@�a7�; �$;�K��pU�@ط�|�ed����R�������U���/�@)��_ƋS�\�1t=El߲$u}�C�闋i�(}}Y�\VV?�����{�)�`I®��AW��}So]͙�Y��I5���ƶ�U���l���˃�Q��!p����o#Yc��L���n_��<v���������E�,�e�1_�J���(3�F,"u���KC��WPj���aa�#���	�� s�kr��>���ik��yS��ypU��v� b�C��V�.g{��<3~Ø�yF8�f T�I��=	wCR�Ձ���P��1=
�D�2�Hz��zc�;���������Y�������݇7� %3VHfR�x@��eC=
㾲=e��n^�2�ԟ�,q2���޳�>�����j��cs BR�ٻ���Ӎ"��rN(���#�$�AƧ�$�jG����ژd$t���?T�,l�?��$�P��cM��/XT�R)sO���+i�J'��k���Z�����?�p�>ya�7#g~Xp�w(������F���Q��un-��;ܩ�dƏcf�;�<DzDWU���
_>��o�+	���+Mp��Y���>a(e�/7�$��T��Y�#�}v2���2���;O��G�d�zW�F�܏�������݇t�@��Sl�5���m$� B*^�a*dg�hFj�l�A�Y�u���d��Λ�p ���]PH����ֽ�iX�Z�RDfa�+�SH�~�$].�<��a���!d�xM�W���/��C�ic<�V�����L2x^Rh0=Ј�r��!;���Ж�B�蕦��:�H=RME[��)�H�$`��|���Hͪힿs�Z>a�`5�nS�0i��I��� BO@
�m�@�a����Ђ^Ҿj#��=X����iv?��'��0d���3������v����R�n̿3N���}�=��?i��+z\{n�������Z�G��Fm&��a 5q+C(/m���2 �B��Kݱ�>���,�Ȩ\�l��B�ŏ�ZN�~�3�z�A�Z����~����M��=�$�4�ЦZ�R�2zs��&�1��>�C{����r���z����Y#}�-r�=N3��@C��T"f�H�*Ӌl(�s��T�q� 'nMxp`Rb�����|��0c���wů���4"5=���=��kE4�̅z�v��R���΍J+�
��9��n�Ř{Ϸ|��n�䒺�-��p��<��w���6b	�,!1�����C.��Ԡ�R�O�i��O�ݪ;%�f�s֤�)�?,	�V�j:m�����z��1G
���1/�>單_=�y�����*SZ� ��&��u��q��ɯD1�AV6�g�ȓIW�q�t�l6�f`��qS&�,��f��cu�+N1��@s\��/�x�l�d)�+؟�C��v^�Ε�8�u��8�O#��Ʈ�x@� )�y��X��w?��"�"��� ����