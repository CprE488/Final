XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�)��`E���ZL�l���g�r+;�C�[]f��s!W[D��t��$d�j��4ܳ��1b~�q�9Tk5rr��%��E|6���$��I}X���B��t���-�����lHѥK��tj����cgU�u!�i��ޔ�'ǐ�#�J���<��9*�2:���gu�6Q��E�℅��
�O��̫7�ąe�5��o�LW\%	&���U��j���O�����;l��'P���l�
�)-�ky��Z�o'x�������1��EQ�8����9��'&|m2b������q��i��6��.�U��$ю��,@G��aۊ�zN��S��ݧ/!dв~�Άq� >GV��� �o���"��h�\�C��6ݹI�ʏF�:H�������K�m�����T��JLtu���ݤ��1�����=_�r���-�Iе\{U������F�������+'������ڃ^�P�/C�������A`�)EB�"h�7f13�e�����vީ�K�
O�G]z�D8�����P���	L�'��Y�+Ђ>h��0�j<���sD_�e��6g�ϝjq�F��ҳ�j7�\fZ����.�~'Bޮ�cj��=�OI;5�q�X�<��������KV����6S�_��$���`��J� n',�/%���a+�d&l�����K�7jq<.�%�,��	�_H�D�������D|��r`B�3��U�	�U������S1.�����}Ɇ���n鍽()��sXlxVHYEB    3fdc    11607s/f�3���d=QL���l�7y
|M�d�<Ei�u]C��A��ۖ�o緣�0��6|��v�i�T�jނ�>V�,�7�Mݓ��)K�_W�f{�WXT�q�'z�.^�ի�����l]��"�>(M���-�h�V}|�^��?`�!ѐ����ve\�A60c2⣉:����@�'��3��\����TM~�W��GI�ő���#�r�e�K��I�$����j�Hc�E�sp~ Z�>}��f�R�4Q������zn9O ��2�A����P�����
!���{�q��po��_���0�^=��;Ɏ��5,�`0�e&���ވ ��ˌ}@L�	w��	�{�%�#7���7�(4�/�݈ID��Y�� y�x9�<t2i�ΧKYnq����6w�^m��ױQ�U��y}��_ߺL� ;��`��L��v��"Z��]�p7[=���D݀G� ��R������j`��F5���_H�x����P�{d�Żˡ�ζR�nE����INOҞL���Z!^k��@J)�@��P����rZ�_��.{�%AD��&z*%ِzZFFg����j�����E�Oo+�R̥G���>s4?CF_�.��$6�V		��7�����)�es���؛|\�8��������J�($�Y������D}��EQk�F��rΗs5���IsJ�2����C_lO��[��
�U}(4E���
�L�B����8�[�1����c�PZ�C<�}o#�ҝM�M9��Q�q�G��J�J��s��'��u��Ҙ<�� �I@R�S�aV�$���𰭶+/��.��%��n\[��Ѹ��pQ�p��c���9����E=�9�uR*.K8��¢���b蠟.l����4*���2�� -�^q�u�W쮋q�LP�mD�6���E4׽dv0�-�5�-�|�� �t�_ߍ��2�w�Uߏ�2�@���{"-�6#�xr��;>�T5ZKf������8F�:�]��>�Y�c�!�Bc%���"lx�J���s���?��tN���;�?_<y�na�����UuQ��h)�S�lA���[,5���&z����dҍ���-���2W:�����f�v N��X�d`������S��{�@|r��/�tn����e�4��W���^!7餧�=���O\�z�4 �<�J����""څJ����By}z6�H3ڿ�T�S6r�F �I��&��Fb��~�2��u��'s��J��lt?I�ȇH㍕�-�C�D�fʓ�vJH���]��7_7�O��;(#�y����:/����-=�@��] �+h�K��b0|���bS�1:k�XI�i��re�7�(�pz�kXc.��9��@X&��:�@��H��x �ģ%���k8u�h�i�u������l���Ǭ�0�G�������b���z�[��K���r���p�w�_t����%�!q�Y��" �#h	l����ơb�vZ�n^Ɠ��ԏ#�jp.q�t���-���0��pqW����k)ʓ��c��W��-;{w��`dmt�(�R��������OzK����:�,��'Y/ձeL�e=��8m��n�4���i�l�F
��J�,��+��ʫ�KC��sD�n~�� #z�5˗��~��6�d�018��~�P��)(X�
�Y�y�SQ=�AG��E�����hkG�f$�'��@ɚ����Km١ׁa��BG�}z��<���Ukluc�{�f�2�b9�-�o��/):vdx~�z�Q��&M�`H�f��<|U��~i��tT��
��<{�2@N6=M��;���g�Z��1����tC�a�f}!�>a���kG�W��1t�K��������Gj�71�ҀSw+��(�v��B~r%��w7��*��y����yiƒ��m�v�o�������w��&���c/p Oͻs �6/��~�>R'Su�p�xe��#ʊ�� ��Hx�DR2`��(��t]��h�VW�@���w��2AHt�E��go�V����	��}�_0���\ �����wr�0�h�+\�kkESח���H=�xl��$�gu�w��肽 ��������G����N���ƏJ��w�96�!����i>�0پ��j�H!�eCM�u�6���x
��ѯQ��DV��-�8��B�ѱ.�ē-u!v���Fc�'��2���4�r�b`�8^��.	zm�/�;�,���M����UXJՏ����{��"���*�F|�%L�m �o������g��`e�:[YO���|��$�s��.L�ݵ��
qf�F�t�����X @�u���Qg�g/[U�`h�a�N�K��^q��L�a�q�~J��H2�rWq�p��W�o_$�ɜ x2��?�疒�:%�[������%����A8�Q��]��U6S���VO�4�-K����m�qzrf����qս�2m�8�JQ�$]{����}��Q����@��L��t�% i���� �)�zsƠ:k!=)��f�;dC��A.Al�gP�,b�ۍ��kc}ʓ{�r� �p���~{�E�&���к�t�
��v����Q�~3[�-�m�d'Jn�˕Wr��62�^��i�uO(�[�a[��^	�Qzx�P�^��o���եA�z�qΠ:Tl�F's���N����:Cz���>��m�t�Uf����r�@��%@��e�Q4��p���5y|x��F!?�@��k�ʭ	?t9P.V��������7�n�l`u�g[�i������h�i)9�L�а��=U�N{!do�� �,�@Y�,*Ƈ	�>�HX�+Cҷ�&R�yk��?�QMk����x�*2���u]��`�R����F��աPK��+�g�(��bV�X5W��6��J�7��>�B�l�Z����n�x�
�yG�1�D4�1����U�[���c�r|�
��v�I[�`������ڀ!������ �L��lN~X�FNC�(�6u�M�6c�*��W��Jz+ذ�5Щ����jQ֘g6`���KS��1}����g��_-��,�e"a8�9�!iQ����� 	3��k��9�..��w�q��J3)U�Xq�8�g=�!� �Q�{�)��H��$\�ܯ
f�
V�`^,p3�៊;r�O�	8UF�d �D���*"p*:��o_y/Ȫ�J� %~�4���ɀ�jĐ�΄�3���J����3�[��2	����Y���
:�v��	��8<�+&��*�H'�]*�W@�O�	�=�E� ��"�I��^�G'U.�B:����]Z�u֘�7\�6��k��䈌_�*7�))Y�$�B���Xd�ދ����b<z�EL�/�g��Nv���{>��r`�dj7,܀��ma�3�p��{��2'$�a�w�:�m�S�4�� ��u�D�u7�KD�����|k��ތ��(Q�J�Lt%�k��k6��(�b���+o��3ٿ}oY�a9	� ���۩y��� CS.A�9�6g_�um�7d�iC�6ɂd����x(��nk�#Ϣ8��`����tHS�_8��������T�
���;�m�����vq��fv�"�h���D��j���N)6��E�Z�ZD�r����T�<��x�e�fnI�<-���q���.-K&ع�^�s$/�G�n��քX���H�������*9�W�>�7q���X�G���*�����#O��A7�Sx�u�X��!�ގ/�2c4��a)"�9V�op�E��ڛ��B�A{X;�,��m��09�v�^D�.�3�e��r#I������D5��X eG���v�l%ކ����.���*�wZ�{�Z�����{�3��.@��0_���W�����tA�u��'��ZM&�dO�\1/H���Fe��r,<%�|�/]R��H	y�8��[
���0�f~��a.Z��C�P��M�Fm�(fH�AK�D�i��&�:C�-��[�!2���U<�{r�3K�H�͉��~�kU�v��T^|��#���t�\�'\Fy���S)$�"�sЪ2AztHesS�Q�x'��%�����6&%!6=����͔�T@����_<�k�͗��O��x/��O���"H#�!��v=wEwa��[� ���tN8�|��#��t�G��6���	ѥ2="�?͑$���L�#,&i��P.�u}���σX-�r� �4�5�����T�����qt1�a7�3?����3V�9:G��@KQ+�[�B�/����\��H\�Y7�U"��q
���;&E�L�o���
;~��~�b�D)N��5N���m�[��f6�R���L
��q�o5�C��y���5� ۻ�Hϓ��K�X