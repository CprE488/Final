XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�ER���v9�����;@�O��E9�1��Aoc�Q��Ɇ]�o���l��ޢƫB,e/Dq��&������j6~J�qo;�.z�����h(�]݃ң�&GK1tY+�`m�3��*v=q�+ۮ��!��@�0�f��1�]2W5��#Sl@�A�c��-���!�W
v�¶:%6�r��4��B۳*ǜ�z�aoѿ��]D��/oz��H�ͦ�֨�����5q���O��LC�(����BG?q������X�e�����޸�7�h�DQ��� �E����3��/0�z;����t�'9��i�=��gͱ�v�Bl�ew�[;��:�`�=v<Rgt.f�$�Yn
D�\;�9����E^>�r�50�s:��s�2���??x���څfn�A�Wú��|�c�[W�\3-���pxӪL�j	-	�Ts�2����������[E���3d��1����i��\���IR�n��`j?���)i"o_���^�t�}��S����9�������r`{U�Q�ᨤ��%p�ؔ�ej���^��?S�&��]�-�TzOhC�@��H�����,?�RQ`�.K�%iM��}�]��\�W�`��\Z�K(X��f?Z���wm��3pcF�we��e����>��^�t\�Zߩe]�4V�����Qzh�8Ʒ͉M$���5+�����`��ܴ���]�&�R`7��KaS(1��V��i+��kS$�<��~6@Z�jL(�gt|/����,�XlxVHYEB    3b09     f80 �=�Fѓ�ܛ��+%�ճ؛K���.�*���#6���a���]a�C��3�XAН��WOi�A�q�4����|;n?� .Nl�E(/��p5���pt��Z<���%�9���l��r0̉�W�6�V1bM��C���?r	c��V�ʪ��U���㷚2���ѷ;�h[=�P���,k��i�+;���F�dR�C�%��G���Q:��I������q`���А|�9KZ�	�JT���&��̵{$=òM�U����H����;�F��=��ٿ��D�Y�,��x��ΗpqX��gX��N�fR�|��H�"����b�$s�$IQy�P�_��M�AN�jZk�m����Ǫ⓺B�yF�Oc�nP"�|�T���NQ�1��1�� ��*�N��������� �����5V���qO���^�E5�i�5Y(l�B�}�O�ޘݣ��7�8Uj)�/c�'��d�Z��Әu8�;s���/�B,-af�!��5)�K�e��k�)w)7#`��K2>�L���%-#gL��S�O��:����nhPm^p{8*�7=�8��>��'ex����]�3��4k�e��w�Z�ϑ��zu�&W��|�4!+����-�b%C	�uA��{E����!�;��g`���&�����牉�?[�/�z�́�|���ᄞ�>l�u$G� y��댬%����qϳ�A}?�Gf��1_X�A��y�)25#��7A.�!Z��yՔD5jhL�ZAM,�7,���XL&�=�51��l&�;Tq�8���'4��UpHM��}�LK�5���Nl���:��Y�S�[?:����k���}zĘ(�e���4�!�FE��� d��-�&��`�Y�Ѻ3�"����9��|y|/��a�/�qme�փ�(�W�������l�ѡn��_a)j?N�fA� }�ר: yO�e�#c"~zn�f��rq���$MD'l~�R�0�R��+�fZ];��هn�jve$�,�]$���[�rP]Z��x�r�4�7��J4|�1~*�iEw&���.�\��� ���zd)���&��`�o_�6�7j�h��%���e�H��m@Й�uW^5�5���j3��E0n �Ǘ��g��f��/p����5�8�	��M!C�j�T�_��(���B�.�u��Z���=����U��x��Yg@����c����:����I�+#m�C^`@��pY����˴ぼ��Q��hNRV��k��#D����|f�u��U*U����q�yQ"�� �R���Z:w_�D�Q+�*��q�/�<��_�۬�w��Iv�Ω���+%8#��ee6nue璤�9��^Э�WfY���j�q.�;.|l̂c���x��4�z+�D����mX����a�@+b]͘"���d�)���������&p��9嘞HA��p�{�j��|��>8iWpL�G�ԾZaZ?Dx*dGK���e\j��T~�zY6�@�77ɣ[% �x�1|�徖�z����qҏ� ��J�a�$c%���C��W��̠����ܵx{l釡>����v�|����\l�q�1Fu���*Ie��[��o`��l�������=�z!�g�en�j�½��������&f���*p�Yk=��:С�c���n�|o"7h�Ţ�����eE��òz9�0�e�2�\�:H��a=�!�fU��o��b}H`���#�bh';�o��Ë��z�EKTbR"�.�_��GQK0�C�b։����˦�w����I���Ӓ�D�Ë�Oi�=f������bx�V���G�r��^0��.75qե<+��m��W>[�նX{I�1xc}�q���c�>6�#�S��E�\�/��_�BQi/R�4T�'źS�b�C����7z.e:������ؐ9vt^an/��_�jg?_�P�i]�ґU�!.i���m�T�JXҏC��jFmpUԨ���W��k��p�[K("��,<��X8?F��C��y�z�.��'��>��x�X�'�DN���u=O�p�K����}��8���a�����d�`��%(��aA���k'��xB�����$R��^s<ss��wy���r�h���mT�	���N��O~���ɒr�����h�]�	Z�2p" ��o1��̂ �o�w ��ʽ@�F��kd%�Ҝ
a�3<��%�>��R�_��v�"���fL�
��D��ܟ���cѐ�����r_���~�53�G!A9}Jo��S^@��q
h��<����PHu��.fL��o�b�R)N�^d�a��,�E�%^܀�ԇ�sD�����?%���-0��b��U�o����������NU_�����.4��b.�<�w}��-�1W�����������C�����<�@~ �b��j5hpn,QҠ0S�=Nc�@}�琬��$��T�u�Y�f��jg� r;�n�����7�l�,�f,z�K�����xQ
��E�U����7L�X
��j���{��v�SRX� �W������]�A�İ��7f2^�@�9Z/�Vk�Dc�󇱃|V�ܢPy�5~5c�t=����l�sJfB~����K���ɗ�U����(ê���B�sV2���<�`f��l�O������x�6�ilz�G�8���/dF�@��V?q��:�ټ��Q'�V66�o
�_��;��~bװ~�L�����P�V��׷,�[!'�#�p��E�0���yD�*ضiƚ�1)r*|>�~'���=��׫P�p=ϐ�
��H�/�#���j��Ň��� F����m�گ���r�������t����p����7���Z�U���| ��.�&E��L�2�}���[�#};���F�����YԴ��1��r�Y���a���d��}�l!��ӌ��[B��+͎D�r��#Iv��ԑ�<�f'G)�=2����h�!�RT��D?)<3��&�R��l�w��Z5�@޸�4���Ьx�p2´5�u�-��݂�X������S-iB���s�����|�:�Y<M[���Xv,n�9�E�[�O�mVU��)S�F��	rW�r����d�ʼ���r�YJ��N�%�$�=G54�V��p�x���Q���I������<�a��_6T��{\~N�'�D�%�@Kl����uh��(e����{q*/��s�n���Q� a��U�
aeM�$�e�����,Rn�Ԕ��/���}�!'5i{q��i(l��:C��7�/2wS��j�]�ΌZ��gna�Jg?���ƏN㩱m��{b�M�����ɨ�'�q��8�ťҰ�	��A��=菏<��-4#(M�e��0kf=;����'�	GZ?���pάedm#��k��Ro/���h�S�O���q��jN���H�8��;K��3%�ׅ��I��+U�`��Y�6e�0���]1"("n0o��*ӸiJ�W���fV�	���ߝ�1�f�3��(k70�S
�{C��C� (W/�ٟ��O�dbP 4%���"g���K,'jy���������h{G�竢?��«��@.Ěӌ��v��k���,��$�}{�ԕ3��!x,:�+!E)ꩅ�� �!P�5�9�sz�wP�D��O�nh%�)�L�׾Έ�RϚ�h�:��P�DО�E�)���=��O3�_��}��k%�R�&����M����� ��D�ٔ���z)���;oeu� ��W�<����B�p�aY�+H	�dg�V,}���yHq�d	���'+6�/�d6��BwB���j'�n��,�- �	��
,���i�ݨ���R��"Q,�R��k��>�D�z����[���]j��M����@��"��g�M������^�\'�4�5B6��