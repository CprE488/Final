XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��t���ҩ��D�A��m��p-��4Z�+Ry�*�\$�J���LA�@�܋�/~uW��m���i�1/�S)�/p=�ۙY�����x��+�(�}Pg�\��&�S\&�=��/�4˴V��:d�N3aʁ(p���&�����/�WK�z2�վr2Yp�-*-Y,�Բ��� ��X�ÂG�;�ְppž\�� ^r�R����p�_�� �d��\�-"��WV8���V��d�m�7�	�9~X���lP�������D6/�tppG��R�8�Rc�k��F�m���z�z�ֶU9���4C6��k��1O�!�6M7XG9T�]e|�n���/�1�i��C/s��'ń�7@����D���5WOX�g`�N|)�?�(ZH͂U'l�������Պ��E!m��1�3?�Jk��IQ�3~ސ���u�˿V&��Z�؛,���$����M�����M�l_���,t@�a���t��ok�R�V�àѬ�>�Uq�=-�5���v}����� NS^��6�T�ԑ�ftG� �e��X=�#�����w3���z��Tg��lUv�7��~^�b��U����y���W���Q��W\��*z'�Ӏa�<ֿ��hv�xL�E�q-�H�)����0֫�(�g@Q�6���\ ��@�xv/E�Y4��ḳ����QM��	}9��۱���r���ō���M�w�m��\�{햧
�Q�0�H+���mi1K_��<����[><���KWq:���3���N�ΟKXlxVHYEB    fa00    2040�u�A �"��=�}*��nZ�NI�`?O�����Jݘfc5�+Ct�%Q{�J����v&Nr�k��uay���ʭ`O��1?�|D�S\���	cV���UIG�	{�4J��`��A���dl��0��&�X���a����5������F�Y�e	?d�.A�By\��N�3�N햜}�5��Z�UG�x�0�D�}��m�^�^DɭL+�̘�)�������X6�B�,���Ly���kƝ���N��ncɪ���8ԫ������;r�����\�s�P����?Q�J繥�D~,�eX��l@��3ޭ^�T$*=��ȭ/�AuaMC������4=�
���U�������̡���to����`�fE�"#��7���C��z�_)v^s�!`��u�|UABB�k�����{�~S{���	�8ɭy#5F	a�][08��es|���ω���w\�����W)+���x<����:�⁼�uΤ<��^�����/�_Bѳ�J�w B��|���������w����3A�z��}/R�����lsE�S�x�e%1�:"q W"bI���aO���C4&M�MbK�`:vz�9��䣥�,�Q�����gD'���b��TP��B0�^�h�H7ub3�BxL�F������%��ޱ%p�/�q�w}�t^�T�B �rI�фh�1|oY���Ϭ�O�٫� 
Z���Q{x>b�xFo9Z��������Z� i$\�V�1�浝����H����@��s��D4[(��y0�K�H���m0�5�Z�����������ܔ>�?:�$~L�]�>r~��}#�|�W� -���'���)+�d(Qa��z�}��«~�c�v��h"<�υs�r�eZ�.it���祀=t���
�٩�4U��5���sȞxΆq#���Ԋ���a�+�'��?߇�Vg�-'�:�ZV�`g#��H���,�������qN Y^L�)�?
N�!�x���dP1� '�����:�<��0b�c�*
v�NC3�xv �Κ���ʅM��1X�?yI"����>5�ܸ4���@F�թ�D�}#s8�������-(�2X&,ɡ�Z����NMc%�Мz����s��8꧈MG��n)���+�UF +#CC��w���_
�y��A���N<7|���K¡^���/���~AӚ�F�Ŝ��'w᣹"���@��En���
Q��+���/�{�2M֚ܖ����(hs�j�� `3;�~ k?U�2A�Zr<��
N����%\�pO�O�|=,���7��O��D���m?�vqD��V���xGJ!�\�M4�5�-�/��8^��,r0?*�7�f�";谻3m���*�g��N�(�gB�3�FR��P�p"��a����۫U�lNn�{�ȶk�D�!�/�]h�wXIWkD���R����\�j/^;�+!�����23el�Q��KcEd�N-������^:vv%Yx�hN��'�.�6�5�<r�tX4���yu���o��S�ğ�N�˝����Gd(j|�?�B��M���Ж�T�ت����	��JM��W��a��	��S�J�����j%ֽ�聋�P0���@�ND8����������[�#����o�Ӈ�����@�Sܰ������n&�$���	�D�[�j
�b��<�Y>��~�E22%�]hH�Fq{��=�&3��ĵ��(��>�Lu��Nbjy�J���O<�ŀ%z�;����f��j;呪T6?r�q*��v���q�p<�Ç��
oCf��oI�#1BB�'��a��h�� ���/xދnq����/���a� BNx"Y89��y$��Vo���pG�V����k����������F��s��h�fj���"}��l�'2ZLw��k�Ik#9Ak�F�Rgډ���&�d��g Żd�`�\w.�Da4-H�$<t����Y .f�w���&^J,���T�V�b#A�SK��%h��E�M�%ឝ��!䆜=�m��r���=���ט�8T<�U�~��;���Ām ����CX�� ,�:��Տp�S�Ѽ����sn��ԓ��H��2�(�v %ʄT1 {5�6�����Zf��V���=���TAk2�n�3�P<�rdP�$M�.��10w��_z�.�Q@[?�}��j�C]���aC�=����ΥD�3���DR����+MH�:+!�Lwv|�V�4i�*�y]�L�(p�eY�&�T�Ɍ��z�y&	*bh������;��1�MW#�� ?�ɿ7�ƱZ͚L�V��[�B/���x�j�爂�����$	����Vt�N݁���>��!���1!J�8r��*�}�6e��`�����ݗZ�[�{�Ð�^}�3����+��$�=�d�mE�����Ol��N�֥
�m{'G����7�p��kM��L��?���3�̦���o�ވHL��*�:���5��2QK<� *�E��D�7����N&�<��N{N'���)͎�]s'8E&,���qN�K�/�$�FC3���ي�O��6���N���5�H-�/	�J ��W�O�E\žB�f����|J(/��*�a�@��(h�w
mM�9s����5f�����)k���և�����h��-�*�["�Nt�,�R���l�U9���k\QW������!�<D:�@M���v5�*�sT�}�tr����fт\�6�Co�jt�d���9�Hұ8Vֹ�����J�γ �'9�4ȗ8.�w�αG��v�Yd�)K��7�Lɰ�U���}���,���(�t4���Go��Is��o=����-9 l1��p&v�$*3���lq��+}���1���W6�q�uRJ�(Tq%�5k�1M�	Tư�9�3�������5𗀭�r.;��tb�XV�F����W����@K�1����C��^輥�ٶ�W��.4����x�Gz,����W4�ʤ��SPD[�.o��)��E��.L���%H.SBC��cV[�]�!b��^{)��>VHO-:j#�G46�E�W��;5���cʮDr�=����s���*� � ���	���\����i�2#w������~VA�)���r#Z��B�/�Ř�(n
���W>���5V�D4�80V���޿F��zx������,�|�?:��S��f����:S�ߵ�cYK���C� 
BX��1���Z�A��^pc2��<LmZ����s5V[ME���B	��廊��ɑ?Z����ϭC�F�i߳���WF�w�����Q$�<k3x��2�P9��u��Pf��:!��l;:�ih��a-l�ک�e3bZOEp����H�_:�o��2�#&f>�O��lP�&�\�Y��A�{�|t���sq������(�o����~$дIN|5�▾�qp�k��LA&~G�g�hC'����;$@2�`�bÁ�M��k�]�ɠ-��&�/ۡ6�#��[���tR�/��"�N����l&ڪH��V_,�AU��O��F�������k�e��U6�%$��N��i^��;������h|B�5o�͙��&1�$gx�p��+���d� ��s��������b[mv�D��a^EX��ʩ����x�)w����ŲQr�VI��%q��.�(њ�����t���}����DQY���z6�w{7��"x�E�v��8.է�/��9:�X�cg�f��Y�zm?��VR�8��L1�zܤ�o3�gj�pW�~��	ߣ_=*+��8�a0#/����!�b�O6ܢ��%�9�cn9�s�C�QF�t�T��\t�?j!��7�ʟ��E�������X&���}3�_ߑb�Y!����1�ݶ)_�dlX�	{�&r�W�3Z8�M��ą���\#�Eώ�	e�$K}Y|oQ�#M�J�,�S,T�RJ�����R� !�W[K!��M@
�zo����@�����.�U��*#&" �����OW(6&�B���'H�?��84�J�^�W1f������LXT��yҨG�n�'vCZ`�r{��&r"`�ίgг/��=3ހ9(���\�o-��I�!lV���DuO�ýBա_�
*�0r:��)�1)8[^$Oz�h&���B��Гz�mTt����Rk��̘�xd'������XY̿.��_{�N�}�O��h����L�=\�X���)���MF&�pM�2o�`|���/z�+���m/�tQ=�����D�z�<ۅ�����mHm�Z��0bв.Y�>K�G藈�E�����5�C\�`�^+`�������D����Z�v]!W|T%h�/.���w
^|�_�N-+��)���L8���\�
+���,�\���thw�t��\�r��F��l�D�$�w���*�]���T��Zj��q`��'uſ��K����\�<(~���.u��R*G
7|Mώ<�}���:iޱjG����Ǥ�J���Q��L9�]���
i� d��V����,f
��&^�k��ŷT3�^yk� ����C�;��� ���6Un�QLd�ƻ��<c�ҥ4�%���%*̋�kd&Z7�7�WgI��� e�U�8��r?�ߢ��6��xV�>ǄѲ�o��=j� wV�4C�J���4�e�5�<zB^�ԡ +�	�6�����W��Γ܋m���P����R�񐔓�q.R`I4�s�F洛��k�j�s7�ϓ��f�;��;�G:h$�����Sl�%$ ����\��C�x��,�������}Oi�)�G�F�>�4i�?��Px3ۭ�s��#j���,��q=	��g�E�+(.)D+	V���)S7���(����̓��dop�Ҳ�.5̢��&�y1A,����c+Ȯ)a3��{��������[/�,Q�-�����6�������,����ot�'�@E�]a�}:ߓ�K�j�]��]S|�q6y��>PM?�U\�P����	��L�*L
T$ʡ�(��XuS���$�����Te��:b?�mX��+ �p�rz�.i��{�U>����T��@w�	��v�;�ڃ���~¤�͖ʦ?&��f���;cAiٲ�G��C�mA���x�"��λʀ_P_��,@������A��Ηzv�N&����Y�����u�jk{�0b[H�=>"  ̦�H����%vºο�`4�?��r/����9�8~KӲ�*(�' ��e��̂+h����L��#����������h8�|�Z?�f�X� ���.K�4ɍh��<=�dhI���S%���#Y������&I�)�H�J���@�Q.T4��h�����)�S"���Y�/�{p �R��/��WV���'�`Ftph�T�����*|�d&�?���:<��!����4�.
!iиސ�>Q��M��=�i�i�soٟ�ҕ�F�Oē@��a���ଓ�vR���}�׉(��BUΎ���W:.�]Bx
ag�\��M"����/�1�T{	�-�UƋ��9�Uɫ#��5b_q��4�<ٗ�+�=�i�����E��s<�_B�i�y�F9�k���b )���H�+\�A��-ô�S�_�8�gaƉ���G/��+\%�}�΍��[��F��rK�sF3�%Γ<�����Ԥ���g�'��w�����2�u��*�Q�Q�g�JӹH�9c9�m�!tjx���,�fѺTF1K��9k����M�\c�)�c�U9~���}*�|O(��WM�֚��fn����+1�:Ʌ��N�1U�W��I:�S���"u/H~�[O6m
a}�w|3�I���=�%����0�^��(�>�6�W]8�٢+�"QxR�6
�;]�\���_̳��t�yr_��ZDBhPV���&�<Rd��)إ�l�h����s�;�DR-�[HW�-ʿt�s���:FS��iS0]�b�Z�t$�f)d�DeO�ef)��y�K|rnq�.)"e�S��s_(Q)o]�����UA�Rp����"�?Υ�8]�.�0�9z3:ؔ\ZL���w��r,8]o��b��	Cl��n����(.��k��`�'���l<����X�2���d�,I��/1cൺdR����-��P|�#&
��9GUdp\e�mń�u��a-� %E�;�u�ݜ����K� '�Gz��U�S1�:�P7�F8�<��l��� i��� �i���o���2t��ox������E���0%�'�^����y�`x��M�������q��v5�` ����,��h��h�"�Z�pk2f����r8���X�[�|���`��H�Ekv'����r8��������=�?�/�A~���8]X�z^��R;��Bh�L�W<��{��cޜK�l:FE)	������4п��H��\��y�Խ7-�m�d�����IQ�Z&;�'���V��	L}��z�����������Ŵ���� �QTO�^%�miI_T�#��E_!&�^���W�X� ����k�8�C�w��I�0G��#�y���ٟ�"֯������jШd�w�6
�#PB����������R�8~�sBØ��/rv��@�:���;�v�y7G9�9@��XpTR�$��BbX��oJ񬝜�0�l���_V�oq y%�n|����ۥ��0����6yb�i��r��Ec��%��ތ{Ո�rĵ�� ��jg@���a	F�����h�[E�vE[n*R�g�����@N)�`�'C�z�+���AfS�!m��E��q{8�WA��/���
v��4g�:������bxX�)���T�N�or��q�j9�ڡxv^!�gã��_����i��%=���J׆���p�|��$U��r< a~�Ȑc6��I�B�e͸�|�4�2㴟�W�0����/G�U�B������K����{5H�/��k*}j&�O����y�����T���(sV^���+JO������u��@��B[� c3�>9�U���O">L��UU�G-�����$KB�#��!d{�������>PJ��S7���%
*w����bE����.�,Pv �JH����bY�����՘��Y���tު+V˽��4l���gY��p�_QbF1S������[�B Tҽ���jAM3�V
��#*?�����C�K1,X����cJ��[!u�(��f��D
�l����=-�?	��gr�]����d��FIk�J��+�%����ݴ�|����6N����g25,���P��.��l�x����B�-��r��*(�:�_�g�c̅�x�/*}�9��~D��ۈ'x� ��Mo�� ���0�Up��l�{}01I�^��l��?w^B�F��G�A�W+?�]��L5�<e2)�B���q?Z�!*���<a'�E�Jq	��.����w��f3���Т��8��X_jEU��O�[0���YXz������V���y��p���`��/k����x� ������o���73��P��IN���\�r�q�'B&銩ym�5ҽ1C*&�JޖT}�O�i$��o/Joj.��v�_'k�Et��D���~E��BY��JTHqr��ݕb;@}@���Q"��M�<�y[$�ϝX�7v��F��z�t���Z*5ݦ�{I�풠3��+:;ʮ ����}����.�v&R�<���y�,Oc�����NW���8b��l��݊\�:�4���\��(�櫻W溕w���o���d,畵O�n����bg�'ptV-�2��*Y�au
�� Y��!��J��-�����(:��j��<K�i�����X��O}���/��Y	nZ����;�5���(ڳQr�%��a�z'��_�*�d���+էx�)YB�܇�*%�75d���$^��[y1@ρ,ꍶ�bP=S�:YB��)���0��Ϛ�͊�ʅHJx,y<r%�:��s�=Y�>�U����r	Y�0#�B1@s�	5q�b�%V۪HӱR�����%O�vLHK��j���^k͌�������b��sc������A����ۧW7�h�Ġ���
�XlxVHYEB    4f62     b50h����_U����	����,���!&���X��ġ�STu�^k!�'ٕ0�캫h8�w
"��2�Wn�\�E!���!'�6YEfY�2l�ưC?��>����ў��Ģ�#SuS�����|Va6ۛ���OU��6��b��=�Yu-�m(�{�y�s�dl���(ypY��T|��T:�y��T���C+*�a�!��
Lk����o4�ngU��y���t;�#��w��M�Kyh&l�^�#v��9 >u0��9w����W��3�E�xN(5
�~6�N��w��h3!;��v�i%E	��L��;�R>�k��8A� ����rZv��h��7�>s���9&�4���9���������	��<ŝW����:�P�*x��{��B	Bb~���ܰ.ݨ��� �W]�(�J���_��_�z���@�aYQ�:�3��'4֞�b�?���PC�3�B�*>cq�G�'���SOFr�=�}��iz�m\�(P�T����6���Y��TV�MA���qq��A�d,H�}��ȸ2�'Ŀ�D�)X~���H � q
�0�ϋ)���:�����h�Sj3'm|�vD�`i�~�=�������ǜy�ž�k
D3��!�paL��o� �����O��u¼H?�u�ϓ'7cxZQ�T1�&(���@͕�tMѮ�a��6( �f,��TyF_v,s������)b�;��B;lCp鄞���#�E��6R�GFw�n0��(i�s����3ZO§��~#�k��j>����)i^H3�^%T_S0̟� s��Z�7����>���P�y{FO��A�zZ$Y�n@��Pn�d����ş�5�U�������u	x�c�L}@�5b��yj��y��e�bL���Ch�R�h�rE���K�X�r�r��Sń�mw����ZFyz��ˠ��-?!�?���:>?N5��Y����#�<E���'�sd���M��2�
2�+(�g����1Y3��X�!�j��δU�G5����z�nhq疗<����o�;���g�4r��b͛����f��&`�;=Z�|~Y��P���I,~i�
n{�CV�Q��v!����!4��}�%�����L�A�_�@�EAI��|�R G_=��A&&f�]����$!\�\ȣ�����mb�Kً`�CB��ʥ�����ɳy!Ρ��ŕ6����t�l�����X[���I#�t9���Ѧ��#��_�d<(`wK��R��"���^�����IԡD����m�����-~�o;Ը���6��4y�Quee&��$o����{��ٔ��Q���xUgA})� |,�)|1ު��ء+�7�m��,��l-��B�K�@Z[����-X�'����Up�Ə��}W#�c��p)��h��?;�����o�[��u>����+���3�������F�ۣ�}�AJ�׭vׯ�׆n�d�s�ʸ��A�����FF�O��V�$�0����"�ӑ�q9� ��C���y�=-V�^��T;��e,��*��5��_e6��M�f��c��F����[��:4�8�����D��G�F�����Ĵ~&=V��Q�?]U��#��n��7f�,��>�A���ڑ4s<e{V����ٖ�z�{��B,�y�9�I�?>��KY��rB��Bl{?�R���6;w.]�!w�M��7��? �'��^����x�u]�g����h�	;�|�V�Z�w��tT9L��çG�Ԓg����@�]�=^���x!x��D��u��
�ݻ�c1�i�y˿'��$��� IB�\��"��vd���ol�	���x8F�-|Tx=QA�	��q��/l�/�v���5��mo��[ߓ�7���eK�A��2(A�u=�mc����?w#g�?�M2�nZ�w"J��)@��9�h�~�-�|w�K�U=4��n��l�߭8��r�IZd_�W�/��(�sv�'��}J�z�� B�qEc���D�jXP��m��<�o8��X~��T@��7y�����>�%�Qxq�A0$��QR���l����SҪ�m��\���B�b�qHѴt^��+��d��-׌t�soD��4���kCC��$���i�!$�{���pG�\������|�Ch
:��Ѵ���ݫ�A��d�*i��	ƱmE�7X���:��#�t����6h�����]d���jtS�[͌���j��$m̓��}�gZ���S K�j��	8�������_�5D�I����<oM���Rl�"�c��hd��o��~�����
����o�R��Oe���s����}�#e�@ޕ��J�}+�`�&Lϳm,Ǜt���4w�ۮ�;����8FP�?g}z��h�����O	�*�Oaq����D��A	�uk}Z6�� @�
�-�I�Yw����GڰU3KsX���.;H��@�x҅2��1�$!�Z�Y�z��6h�i ��i�!�b����7f�?�쀷��"�K����$E�S5���;!ė�h5���%]<�-W)�����D҉Wo:be,s�sׂ����i&���8]��Hp�����8֥MB�~�J3��U�Z�#u?S  G��G�t�N\Z`�E����"a�눤#X�Og��O��O(���L(Gm�k����Qo���fU	M�-m���h��O�T����"�#�j&�i#%��T�wn���	��Vl���tu˸�T"���۞zު,U��o��(�fof����>��b�}Xyo#5���\�>�Ϟ�}ӳfp����	{lC��6�E$�t=� y�Z��8 �@z�_]d%Sze1}1.-�ĕ�-�[[�W(JOp?�t�U�H��f�