XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��lr�@��nr��@;Q��<��ф�K��"�!�i�F7{���n��PN��������-H��1���rIR���V�c��yw[U�����ڕZ�[b�b�E����u$�M���^G���[g_��ծ�`P>ݰ��}i�,�A�{�X����z�M[�̲k.kb�Hx��۽3���T�	��v1.���E�V��H�(Ns^��i�G9���K�N�D��ˆ����������B�촬`�}�_�U�}�t��	�sU�R�Bh�Pie�|��1�����F��ZL:M�]��$��Ɣ�'*˷�s�.'���sA��;@��-U+�N�������"͛u����B��?���o��POh
V�t��1tĳ��HT�� Urﴸ!�G��*	FaI��H�A�6�F|P�v>�Vl�c�β�˘B�k�6�� �*�~�~a6�c���9�W��OyE�_Ix����Ve в6����Z��nG�N�_�n4��.��:2�)55��n�7��W�$��i �<����*K���-��e"��6�ãF|R�B��h��^�	�Y:�T�-��Iw\H{�`�H�v��p�T'���.��sR�-�*d(���I��\.��Z�v����*���/y8a���=/�������G 0�Ș琍 lKv���M��u�U���c���	�?��b'�P+P�h�c�8B���w7���@a`E=�p��`�~��pB���?�@{�=XlxVHYEB    6014    1840%�m��V��}��Xx7�eDv?���^�i�6���}7�nx.���||'�ԱA9�G{���u�=�ӄ�Ɇ�`�k�d��N��'�=Vj���?��E�@���\=#�.��Z%����V���<boxK�%��\㔕NϑP��i�i��<�%xD�t&&ַO��_�����>�Ck��s�Z�	t>�Y="ry� �[�>�k��_	j�}aI_��|ԝôSX�>�Z�K�upu@��ءv�Zj�۽E� �&�9y�Y_U����s���KcծK��0�7��(��@������4O�[_ف��u/�Ɵ5�Q�����Ř�}�(���ɨi�G5�>��u�h�La�$�C6����|r��B�%��Հ
\*��BN��`傰���U�i�^�B��PI�C�~t��>v>~6�:�N?}��x=�r����61���H.>!��q�~�2�"���[��|r����s'�d}M��0��O,Ѧ��{�B�B���31����,ɭ��!�h?�`��嗙^&w�6�Vm
����X�a�La�Op!���'�����&`K�����t��%*�G���)Հ�I5�	4O�F�����<�8P��	z��}�a�0���U�0��O%ϵ�l�-r ��ڮ����߮�h�G��0o��P��v�����!���EJ��C�h��Nc2K�O������ԣ��� ��]X�K�����$G��t�[��L�%��ǂ�`N{ �ͬ"����N���9�#0D��# ]�@��3/V�K���"ޖf �[������o��x�
��9����STN#�B�� �Z�	923 R�
LۙnP��x�Z�3�b��u<���z1v�e�!��dc}o��[�1OR��b8��,������ܓ�Y@���!���K�7w:u���3�75�-�����Du6Ľ�����8����+���ȳV�i�_w�o�k��O��_����6��I��I��|+��Mu�y�6(�[�E�4�'��q����J�6�����؁0|u	����3Z֕��u��t��������~�N~6�f��^0�?� �n��Yՠǌ~�/�$�?"<�w��˩�	�~мɩs�Q&��%j�M���Ax䙾�(������|7JA.!�1Q���܎�~� ���D�<�hZ�1��L���r�~��L�O��#b �$��g�<G�h7���U�rd����[F)�t��!�/�)�J�R�|<��6,��j�}*$�<ND����/��a	P{z<T��J�ǲby]%4OC��4E�����0����!��_{���C�	Y�5@d���P�����S'��/WvP���Fl5�m� k>��G���++�+�M ��� � �~s��K@�����D��u3������p��r8��ee�5?9Ka����fԱ�[n����x	vN���l5J��n`����5�*��n���ti��%���ƙ"�!f2�M��"��w���(�38��
8���	H���[�*.24�۬P���9�@�������e�PE�|'�3�p����D�u��y4��;�=wt	��c����+i����6qt:������~^0����$>�?��w��B���΢��� �������N������h���Z��0A6�ą�k9OJ�u�؁��ڄ�H�D�"�MG�y?�
C�}��u������W�M8½�NM;�:��a����A��5�G�ܣ\��A�d_���}�.��Et@�����������B�.����O���PŐӢgb`ё��	�]{NX��!����5�tY��`d�����Q�k00.�*����3�ƌ��97L��No�Yc�jlŊI�9��,��!ժ�����+l�Q��(��w$|4��\�w��e��Oα{cg��J���!j�*@m�z���=���v{#���rP{��MO�ʖ�u,ǵ�����V.a��� "6��e��e�v�De�~#�>�7R�t��J�-���[���dK!��T���/#�}��M�$3�1M�!��� �a ��ߚ)׽�Gg�`2�16A�O��O�sH��J՜��Iq&�ҝwk��^~9Xol�x���� љӔըTL�?������a���������AUw��/���yl��(8�e�]��D>���m*��A���N�]�]�rC�ΊC�������	`7_�����u�����0_.wt8r㴁-��ع���G�����R7��Ǡ��y��'^MZ{q�J��U#w�5eX�PG����S�1�G�,��9�(1�w-4=V�z�4�q@��]��z^~T�Oo����?�R��eu��;<:���������=(w����5mW�����i�:Sc��K��d�f,sp*Szb͋ZXX���pNYptڎ���	P�_�f�o�%�Nk
'_��B�t�}�����{_�#�^�;����Ua|]Qv��	bRz�{��������a���fe��G�i"�*eP#�����J?l(�����f�ǉ��f��^�/_T���mW�v��j���_=sib�A�O�
���K��4*������4Q�}�>�o<`�[�|6�o���,i��u�)N @�C�b�J��C�e����8�Ѡ�����c��j 9��*��A� ��������z���z��ֹ�R�A+��"7�����!��6��O�O��YƓ�`�T��&�d�ؑ>P�C��,$��k���jP]��_�ѥ2L�` �4�󙪠[Hy�r?4ɭw/ʶ�o	]�^�yK���=�� � ��Isٳ�!��n��\�F��c
��J��Ea2��:8�Wx@���5�@:�tf&��qS1��|�ЕH�La��Ǘ3O0DK �Ld��)]����Sv`�Uy	+-��8TM��c���U�/���0U�)U�p"z�!�,�)Uy�ZDV�,�B���«ڝ$�4�K�=-�:���A��>��Z5� [�v՚#K�s�I�U�3� K�b�-8�W����gyXf���r�.kV}�`K{�$3&�&���<۾Dyr�.�_rC�-�	��ayAT���;u�_J��q�<����~�)��{tQ�X�_�iLm�#���+gqv`������@<3u���2\��η���B�aH�Q���Z$��v4���룼��/�q��?��\��5���.[j�d�.Y��CYj�4�enS��3��e���k���j�5�$1�/j��.3ك�{���@_)��Av�"׃R�\u��U)'��{Y?�`O��]��*ʹ����}G�F�eW{�h� �{#֮tS��K��D�
y�<Ǖ�����U�[t�P�=�!ٔ(�zV���{!Es��_��r�-]x���c��<�\���"�Y���t�l�����|�|��y��o\��Ͻ����q��1c�� ��NGv=�x3}��F87��g 9[�o|=��8M�	a����e�����\���Y��o��(>����o���bh�Sov��DX��5�]b��}@��/qkMM�>�1���u�ʦ����sl�P�DK�J!_���F�G���,WK^�>'~K���X�m�̳ w(.w3�Q/;Y��a��p	-��:��My=�ɣp|�Jn::�?X!AGZE���`���B�7>vds*Hy&C��e�JV����D���b��	QD�8۴p�ja�뙹�s܆�O�x�U����z!�Fۺv�	�s�W��ز���],�9)�M�Dv%�¨9}+�dF�m�X��"��,ƋKD%���16ѻ��Z�	d@���$�9��}1׀��<;E��]�����}BSb���U��$��@��-����[��]g;�q���>Z������C��J����B����f,q��&<�W��k�j�A�OB����2Z��*�'��}�ҝ�i�<�s@�pӊZ��in���� �7��)d��}V�ߡ1�OC��Gr���-؇�I��t�r���^M��Kn�W6�k	���V�p��^i��g�&}��%x��~fz��R��N�_}�)���E���US\�\�9�Qd�M`�-�r�x�
�Y�l��Η�����<vu����_���>CB�a=Q�R����wЕz�L|F�-HPb�X���:�>=@�C.�ΨCv�~����a`�L��uD45���"���'�������6�ل�k_g:��0����6���Q!�	����;810;�GT�$�.�{&�w�Pl��v���M*c�f�\���Ax�q�\��ZN/E��vtpE��;�$���:[�R��PDR�+�|�֞��]'��w8�(����ĥj�dũ��q\�F`|�X%��linf	�L�&"{��({և�c��kt��39`����K�P��0Lʮp���#��!H�,��[��k	�y��脃�]^r��(Ü�4���N���ÿ����q��n ��Ş�����李�) �[�o�VIO��hL�z!G��l�E�}.�(��TL�0i�����F��6I���r�/g<hA��J1)x?pŒ�d�1I�8�&��;�aٓk�ի\�N)݇�f\Aȴ;B�,��`�܅Z��*	Ø*=��8�|̉b���mGҚ	g�Xĩ��+�~0�=��i�|c��}:h!m����5Y�o��M�����sVG���C�6�Ʊ�mb�e�/E����=n���7�*�ʜ�4���틥�+{Te������e���sQ���4���nĮ�\הp4��[�631A}4�+zf��0�����L������[��y(�Z����x�`F����w*�LX$��.�[u �Λ	*{�sN�+8SA��y�s��b9O��<��d�U��U�B�\Օ��d84�++�[W�$��t^S?뢛��[�߇�C���2v�3���N���(�){�է���a��#�y��4_X�|0i�e[ώ�sY=s�0��i�	3��Vb9������A������D�?s����X�䡘v�ƚ�va?��n𢻩Yt�N_�`�3z6�i]�F�3����j�*�\Ѻ%:A���f���~|CG�!Bk�%p�"�)W�$�ve��ۋ�og�ˡ�Qu��H1b
iGڸް�J�W$�c���;J��X�l�с~�Y���\�G]���-1���n��U�}����ٺ��|$�R�D��9w��xT��a!$�8�O{��3N���]fgK��I/&-9W��PV����Qm�ʇ��k�iWQμ��"K7�q�,TB�ʾ���?���c˕u�����I�x����?�s���(��K-#��<�:��tM�Qkj�à�3�O�e�����m�c>�_���gź���
*R�$���_Q (���l)�M��L�m�����������WwB�\�~Dj���D\�u<o�l�����}���0Z�B��KHu\�^H��Fk��F�<�	TV�h�n�M1 Pi
�%-�#0i�N�N0������7�(8��lL����҅0��ez�n4ϔ�ZXQ��I��vӒ�k�.�o��ݤ��Ar���0좷|u�n�6/�_M#����(��D�mL�3�'�Ca�nF���0tn�q���a5������=��Б��vu��+3��g�ӣ����'9)��-*Lbmd���o�:��tXIϳ�V��ﷲn��9�Um�&�݇=���K�����kKO.�t�wuz�o3��9C�����O��%	���&�ŦUݺ�C;f/�h�����M��(fN��p��g<��Lg5��^�pǴ��g��{	0h/�'��D�;DS��QC'>�>�J�I.��ć��PjN����W��A��~y
�8�-g��E��ۀ�'n��N`)4I:�����;�l��͂L����<���K��?�{�C�`ō2��K+���w�A��-T����%=,B��O�<�.z"��mPߦ�>?n�V�`�&��u�]�ᦺ��3�i���Yu�F��|0��g"���-Z�u���`8_1mK��JH�jS`��k�u@���o�k�ﵖױ��(lЋ�+	��}'W��)o��s��U�������K�_I�4�Q�ׂ�t��#�˴Tbʶ�7�눪��ˁ�(�~2