XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ˁ>q�hҀ|Eh)���B`CS�ĺ����4$���*���i=�¿��cQ5�1N����׺b�!؏5��(o,5H�(^�#������:{tđ+Ň�Y_[<O�|ǁk���؂N�������:�)�ށ�3�aY��.�5�8�O�Ø�AF$�x{�N{�k
4X�--�>b�Jm�Qݏj�0r�wb����g��ӕf!O$.��d�&͋b��'��c�0����/��(p���U��,�Ԗ/c�6M �TS��%&~��Jbm}�� �;ы�f4b��U)]j2�y��as��N��]��A��2���a�/Q��x�����Z��v@Y'����e�[��ã�O�6���I���X�d��V+g��VN�Ktd�n?J�A���n��s]~iT i���7Ԃ�$�B�5��Q>45�#��
�H"��ά�L��&N�n����^��6���Qv��!�S-���2d��YR�Еv�= �/�w�#-�!�I:n��F]��$�p�:�Q�O?_(i�U�[�C���^n�C�JGqYw�*j��6��g�hUosH	����pC�-����HHH��|�Vd�_���z�Y��ru��p+����i�7~9� ���os�6��.���v��f0��c���NK3SZuKw�J��G�3Ѱ�$���k73["�h̉D�
����N+�G5X��Y]��i�ߛ;���w�t�f�;f�`.��l4Tq+Eq����BO��_-Al���	�BZ��d'K�XlxVHYEB    95d3    18d0� P���F�%��t쾛n���[��p�.n�{��k[��Y��cj�8���UN�TM��qoV���Cl�̰ksW�N:&�!�[3W
{�t�n 5�ǋ-�I��[���~n1{�z�qu�&�5}A`>>�:P�1j�rN��)cQ$g�_X��Q'�	IT��KҦ|��9�SS��xs��/�O��a��|m�S�-r�1�(���ʇ����B�q���E!������S�?��7�ɨ#S'�Ȍ�p$oſlV��@� դ��X`}����N����*���u7������$ %)�G��������nU�^�� �ؔ;@�Y��J����������/���{z8RW�W	~~��c�joûC���W:u��A���SO�Ѧ_lL��I�m����[^��T GK�3�B�'[R#��X/��=PX���|�C����� �޶̡~���^~-�A��R�!)Ò�����m����n�1�2V�F�c��)��,��������Ez�c�)_�_q��ucd$��2r���ҌBnO�&��K�A��c �_/��x�L��aˀ���(����*���0�5	���.��q��L��k<*�y�����[71�q�F�]/ �.ꜿH\�w��h��[������-`���1��`7aJ�ʄ|�W�wfe�L@�,yX��r%ӂ�����K�L:��;�#��(ĝ3�[d�Q��==��f��1��?{}�A��K���`?H�	=�O�������8������t���<�8tA}M�6l�N�*>i��ߓ� s���Tw�1���7��"����e�W2������bl�m����������{  +�r��|P�
T?�1ֶ�Y�^_,%t�ߘ�ʷ3?�	o|eϥ@)N���z��_�D�l�H��sa�Wؼb1�RQ9H^r��%r����+ֱ����%� \���-<��i[�B�*���S4Q�mI�ě�\^3fo�/��&�h���}�2�J��ׯ��JÐ�X��CUYNm���h�����y$�b���HtsQ����d�y��צf�18=�M"�4sx�ỉ��*:�NC4n��F��M�4�oR��qج9A�Τ�T?q ;y�|6�w��3J{��Z)[[������&{i�jE�m�7
s`��K���ðe�Ft�X��Hذ-4�G�&w+>* �tX��维>a��D�Bx=A��Q���n��w�VcMN��TR�a�E�I�p��*�S�p/8�E]�Bŀ|�h�CU�������_$||a����O뮲eO��\J>\�!�]�-�+`״��}��o�l����xp�uO�'��'��*����O[g�	���D�E]N�������~�gY?R-�<�������>���Б�@�?E����*@���bh���U�����F��/��ȹ�a�LD���p��F����'�d�5T��y�Bk�9�������=WB���T�������3K�rR�\���H�����
��l����PVᔅ�WL�����cH	�	:��t��Kl�?6,)��_v��]��6	��JU"�aJs<q�hyl�"nޑoi�܎"���8��͗�ϴ�'j�q���*�
�"�:t�`*و�E�Ϣ�M@Va����R����P2+X��/�u_�	5�bBk��{V��*�_�!�`���뎆�&��0[Y��~�Ts� k3��W��܍Lg��羟.�����O�Ѳz�8APn��WaHUF�,���+v��'q�
�3�6�21heF֥��H�-$�q���A��
SLKe���ER�k]r���A�rf%@�+M��7C����H3�*�	�<����X������ۭA�#s}7\y]	5�>�9ݒg-K͔���B��F���t-~W&��]�#5��	S���ں�H,�R�?ͽӶ�_>���F�x�B�Sz����rB��W����J��6�����|.ք٤~�PMv=��#��'.%]y�g�� �k��!���~b����:kF#�g��!��)OI'.���X��4�෻����W\�#�Ch�:�?�N̉01w�x�JcW,�j��z�)��~2�/�0�/�X�DΠ\�G�QR�!�j��t�YfRϷ��fm��9������tp�����5h�e]�^��:��L3Ăj�uE��
����:İ��o���I�jm=#���Hݺ,���6�t2�8t��#�9�����A]	C��@�XY	Ȭ�DyV�tƁD��;\�K�gX��a<�4Wjk.�Yn��ִ���	$t�<�-�S��ORP�l&��|�[�[i��)N=!5�����~)<;n�W��?�{����Xm��i��P��:Uyɾ�� `j�[��R�Lxʠ�9�^5zv�w����!CI_�$�`"&���B �P��e�m:`�`�Ж.���U�,8�Sj�
�ג%�"7��ŋr0��I�m�5��7ٖ����(H��=.SS���c�O�2��%�e�C�!��k�4�4r�������a{m-�y�{�5F��ye�￫���h8�-$N�i�����w79���@w�`��)�B���������>�1�"��.���E�"Q�mK�2�jO���%y��ӆ���'}�r���%�L��z��T�F�g�W��FT�pn�)�:O��WZ��U��'�f����]�]QU�;�W�g��M�c���v����n�
>��	㕖d�l��q�%˶�6� �Vrt���^�ی��O䳽F���,}!PGIi)Rt H�L�tqn�8Po�B��E-����SC����B��FT��eu|G���#?�}��$}�ԂSk��
��&C��7M��9#��>�f����&V
jGV����ᠳ�F�� �0��Ƨ;%U�1�շ��H��l&�����%���N$0��g�J��5���zJ\��������g��xT��p��_�G�9�!�9��f�����ø_J�Z={}�E2����Xvu䓐�=��v����1������.��r[N�5�;f�XG���b��`�AhX$���juH#=�� 1{ms��@�d����!�hì �r��ۚq���Cƾ���.�at#�1�p�C��-�o��4Kf�34>\#�o���)cy������"�(�g���Y|�uI]؅G�= �§��Y4�a��^HOD6(�����{1FS/1�k6��Pۇ�4f�s�Ͷ��\>]���6@=��B^�J,M&�j��i�T�*H,���wˬ���>
^D��p����sT��.�)�[�M��~��6�֕����]�Z��5���{������Y�y�H�}CP�%�{�>0ꬕCG0?r�ڵ��O����,���9��S�Y��|$��`5'�A��8��c,]�5ӘOJ�z��	A�������m���{�(<�?��������r�:S;�P�B�
#�Q�R������5�O�v/��ïy�S�5��R*N��ݖ�] ���5�2���,�>\+:1�@���F4�V��:?JuJ�=�i�j�o�Zv=�F�;8�%?7%T��G!X�2췽��l�<���l��BS�
m��>rh�6����a��%���M�����{����v�*�?qEڛ�-6;Z��3sŐ4C�@�[%$/u�{�,���h���\��0���L��_���3�[�WU>h&}+�k�y�q*+=�6�^0v���T��#2+���@����T��wU�+aKE�/�{7�ۨ�ۆ�G~?��}�-k�p�lR�,�s5S���j�1�26��5��PW���.&�;��z�����R<����X��K�Ì,J����ڟaj��y���(�0$6��d@���՟b��gDAj��� =�Ny0�ݎ��1�1wd�!TX��(�ag��.��3���5����S�ZMu����~�\8��x�pK+�m��x�ts�iZ���3�"f��I����&��1��ݧ[,�M�5��m�$ۀ,�P1��G������s���rK<F'}���/�[UB��PW�)���y(�T�/�!�%���xEw�Q~�}�ۏ:��x%�S�V:�g�u2��*X��n,S]��ɕ\E�h<�4�Q�D0�_TQ-fn��(��5�U��n�Vn6M^JK�8#2,$�φ���K��`q�p��*�LU�v�`d]jXWg��L�kI�8�K�'i��jX�5�2^^?ET0m��u��[�"�e�c%B��lx�Z�q���_�Mh��Omu���]�=e�}��}ae�+�%�Կ��T��!�uw-�z��=&?O�ę�'��ӥ�d���Y�+���^���{�ZD:%MA倪��%Ɯw�o1}l{ts��Ƣ�Ea��S�wJeC͘�E��󍃰p�� ����7L��W�3��Upe���ѓC��t��^��6��r]��a+DstӵC�z���:w0M_��`E�Kşr29��ʧ7�+!���.��2�}R�h/3��᥼F�ᇟ�56y��?7���O�n�r�\8	�V�d�\*:�Іd������ӤKW�Lo��u��4���Ո�^�<i�i�����]�����^�乊m���Ϛ��m����T4��8�����t����c[�t3��ҪuQ���w@ҽ���N����c聵}_{>�^�ar�x�F��E�.�����:^�"h�!�	�׵����A��wiqJj��5����m9;f9Z��\�����u�x:m��`S )L�n�nO��/������(ܽƕxz��bD�� �pu����hX����I�D��!�j��W���̏�-}C��Ij5��k4,���Q% B/��&e����%���$H!w�O�V������G��"ݘ���r%>xd[Z��Ѵ�q����G$i�t������.�YX�nw�8�RA*h��M:�Ze�������iIx���p�L���#�� ��ϼ\n��,�ړ[�6:եp���X�ӿ��F
#�)C\�Uͤ����k͞o_�N��y�@�ӈx��<X�"��1�J�"F`�֓��}�	�V�m��&iZ��'��g����Q���e��N+z��:��<�� <lR��h� ���IB�7���đ~SY�t���83]����{B7���������qP	:;V�ן!�kj��^dVf3�ׅ��e�q���:yp���F�n������`n������M?�xUB��u�A�c�/}�I���[��߯�E�6N���b��o�..f�z� t�~H�iS~r�a�e���L8x���_gd��@�"70�ߧun��P?�\���x�2೪*c��G�$*4�,;Nc�=b���"�n1{�\�ǳ\��A/�.p�@���PmXzs'���{�����り�`T<���;͑	��'V�bìB�(�܋�-BT"��4�u���PY^����K���Z��N���IyR�]�h Cv�'d�ŪX��@������5byAO��)᠎�&�>X�F��@,?-3J�O`))�'���{�;n2mQ耘Ԥ���)��=	j_}��>V�4�zO�L K|0u_[m;=T�J�YB�Y��ԇ�u�Q$ݓ�غq�����dF��mG��#��Ǯn��%����i��A�x�� > y���50z6$��񁳴%:����
+9��]�~l3��y��.�94��MI�F�Q1��]��,�d����rPD�h
��O4_;���)"$��y���/�\\�Z�`N'�2����6Td^��p�K��:���t1f{ԝˇe\F��-�iY��uވ�
��ӥP�V���,��N'"wYlN�ag�Đ�����L��fk� l��FUp�?؂إ�m�h�6�e2�^�^�Aqv1�1:�OK��������C`W������Y���B��E�F����07�:��U%�=�Yy3�)��2��%q�Yo�E���Z��w�/�����X�M��^���l�l���}sF��.L��\�܄�tj,������|����
O�ucze�����4��3���Y��4�a�ٻ���Pø�a�!;��d�Ma��!��n ���b�,��u�¨<q#�D�o�cb�~��ۮ����u�	�p���c�����w +!Xj����*�(�X��D�q��}S8Yi9mS�X#'��^	��Y�ݟ��9��*f��N`��sN������y�Q�U�n��Ȃ�d��q-��=��c`;����